// This is the unpowered netlist.
module wrapped_simon_game (active,
    wb_clk_i,
    io_in,
    io_oeb,
    io_out,
    la1_data_in,
    la1_data_out,
    la1_oenb);
 input active;
 input wb_clk_i;
 input [37:0] io_in;
 inout [37:0] io_oeb;
 inout [37:0] io_out;
 input [31:0] la1_data_in;
 inout [31:0] la1_data_out;
 input [31:0] la1_oenb;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire clknet_0_wb_clk_i;
 wire \simon0.led[0] ;
 wire \simon0.led[1] ;
 wire \simon0.led[2] ;
 wire \simon0.led[3] ;
 wire \simon0.millis_counter[0] ;
 wire \simon0.millis_counter[1] ;
 wire \simon0.millis_counter[2] ;
 wire \simon0.millis_counter[3] ;
 wire \simon0.millis_counter[4] ;
 wire \simon0.millis_counter[5] ;
 wire \simon0.millis_counter[6] ;
 wire \simon0.millis_counter[7] ;
 wire \simon0.millis_counter[8] ;
 wire \simon0.millis_counter[9] ;
 wire \simon0.next_random[0] ;
 wire \simon0.next_random[1] ;
 wire \simon0.play1.freq[0] ;
 wire \simon0.play1.freq[1] ;
 wire \simon0.play1.freq[2] ;
 wire \simon0.play1.freq[3] ;
 wire \simon0.play1.freq[4] ;
 wire \simon0.play1.freq[5] ;
 wire \simon0.play1.freq[6] ;
 wire \simon0.play1.freq[7] ;
 wire \simon0.play1.freq[8] ;
 wire \simon0.play1.freq[9] ;
 wire \simon0.play1.sound ;
 wire \simon0.play1.tick_counter[0] ;
 wire \simon0.play1.tick_counter[10] ;
 wire \simon0.play1.tick_counter[11] ;
 wire \simon0.play1.tick_counter[12] ;
 wire \simon0.play1.tick_counter[13] ;
 wire \simon0.play1.tick_counter[14] ;
 wire \simon0.play1.tick_counter[15] ;
 wire \simon0.play1.tick_counter[16] ;
 wire \simon0.play1.tick_counter[17] ;
 wire \simon0.play1.tick_counter[18] ;
 wire \simon0.play1.tick_counter[19] ;
 wire \simon0.play1.tick_counter[1] ;
 wire \simon0.play1.tick_counter[20] ;
 wire \simon0.play1.tick_counter[21] ;
 wire \simon0.play1.tick_counter[22] ;
 wire \simon0.play1.tick_counter[23] ;
 wire \simon0.play1.tick_counter[24] ;
 wire \simon0.play1.tick_counter[25] ;
 wire \simon0.play1.tick_counter[26] ;
 wire \simon0.play1.tick_counter[27] ;
 wire \simon0.play1.tick_counter[28] ;
 wire \simon0.play1.tick_counter[29] ;
 wire \simon0.play1.tick_counter[2] ;
 wire \simon0.play1.tick_counter[30] ;
 wire \simon0.play1.tick_counter[31] ;
 wire \simon0.play1.tick_counter[3] ;
 wire \simon0.play1.tick_counter[4] ;
 wire \simon0.play1.tick_counter[5] ;
 wire \simon0.play1.tick_counter[6] ;
 wire \simon0.play1.tick_counter[7] ;
 wire \simon0.play1.tick_counter[8] ;
 wire \simon0.play1.tick_counter[9] ;
 wire \simon0.seq[0][0] ;
 wire \simon0.seq[0][1] ;
 wire \simon0.seq[10][0] ;
 wire \simon0.seq[10][1] ;
 wire \simon0.seq[11][0] ;
 wire \simon0.seq[11][1] ;
 wire \simon0.seq[12][0] ;
 wire \simon0.seq[12][1] ;
 wire \simon0.seq[13][0] ;
 wire \simon0.seq[13][1] ;
 wire \simon0.seq[14][0] ;
 wire \simon0.seq[14][1] ;
 wire \simon0.seq[15][0] ;
 wire \simon0.seq[15][1] ;
 wire \simon0.seq[16][0] ;
 wire \simon0.seq[16][1] ;
 wire \simon0.seq[17][0] ;
 wire \simon0.seq[17][1] ;
 wire \simon0.seq[18][0] ;
 wire \simon0.seq[18][1] ;
 wire \simon0.seq[19][0] ;
 wire \simon0.seq[19][1] ;
 wire \simon0.seq[1][0] ;
 wire \simon0.seq[1][1] ;
 wire \simon0.seq[20][0] ;
 wire \simon0.seq[20][1] ;
 wire \simon0.seq[21][0] ;
 wire \simon0.seq[21][1] ;
 wire \simon0.seq[22][0] ;
 wire \simon0.seq[22][1] ;
 wire \simon0.seq[23][0] ;
 wire \simon0.seq[23][1] ;
 wire \simon0.seq[24][0] ;
 wire \simon0.seq[24][1] ;
 wire \simon0.seq[25][0] ;
 wire \simon0.seq[25][1] ;
 wire \simon0.seq[26][0] ;
 wire \simon0.seq[26][1] ;
 wire \simon0.seq[27][0] ;
 wire \simon0.seq[27][1] ;
 wire \simon0.seq[28][0] ;
 wire \simon0.seq[28][1] ;
 wire \simon0.seq[29][0] ;
 wire \simon0.seq[29][1] ;
 wire \simon0.seq[2][0] ;
 wire \simon0.seq[2][1] ;
 wire \simon0.seq[30][0] ;
 wire \simon0.seq[30][1] ;
 wire \simon0.seq[31][0] ;
 wire \simon0.seq[31][1] ;
 wire \simon0.seq[3][0] ;
 wire \simon0.seq[3][1] ;
 wire \simon0.seq[4][0] ;
 wire \simon0.seq[4][1] ;
 wire \simon0.seq[5][0] ;
 wire \simon0.seq[5][1] ;
 wire \simon0.seq[6][0] ;
 wire \simon0.seq[6][1] ;
 wire \simon0.seq[7][0] ;
 wire \simon0.seq[7][1] ;
 wire \simon0.seq[8][0] ;
 wire \simon0.seq[8][1] ;
 wire \simon0.seq[9][0] ;
 wire \simon0.seq[9][1] ;
 wire \simon0.seq_counter[0] ;
 wire \simon0.seq_counter[1] ;
 wire \simon0.seq_counter[2] ;
 wire \simon0.seq_counter[3] ;
 wire \simon0.seq_counter[4] ;
 wire \simon0.seq_length[0] ;
 wire \simon0.seq_length[1] ;
 wire \simon0.seq_length[2] ;
 wire \simon0.seq_length[3] ;
 wire \simon0.seq_length[4] ;
 wire \simon0.state[0] ;
 wire \simon0.state[1] ;
 wire \simon0.state[2] ;
 wire \simon0.state[3] ;
 wire \simon0.state[4] ;
 wire \simon0.state[5] ;
 wire \simon0.state[6] ;
 wire \simon0.state[7] ;
 wire \simon0.tick_counter[0] ;
 wire \simon0.tick_counter[10] ;
 wire \simon0.tick_counter[11] ;
 wire \simon0.tick_counter[12] ;
 wire \simon0.tick_counter[13] ;
 wire \simon0.tick_counter[14] ;
 wire \simon0.tick_counter[15] ;
 wire \simon0.tick_counter[1] ;
 wire \simon0.tick_counter[2] ;
 wire \simon0.tick_counter[3] ;
 wire \simon0.tick_counter[4] ;
 wire \simon0.tick_counter[5] ;
 wire \simon0.tick_counter[6] ;
 wire \simon0.tick_counter[7] ;
 wire \simon0.tick_counter[8] ;
 wire \simon0.tick_counter[9] ;
 wire \simon0.tone_sequence_counter[0] ;
 wire \simon0.tone_sequence_counter[1] ;
 wire \simon0.tone_sequence_counter[2] ;
 wire \simon0.user_input[0] ;
 wire \simon0.user_input[1] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire clknet_4_0_0_wb_clk_i;
 wire clknet_4_1_0_wb_clk_i;
 wire clknet_4_2_0_wb_clk_i;
 wire clknet_4_3_0_wb_clk_i;
 wire clknet_4_4_0_wb_clk_i;
 wire clknet_4_5_0_wb_clk_i;
 wire clknet_4_6_0_wb_clk_i;
 wire clknet_4_7_0_wb_clk_i;
 wire clknet_4_8_0_wb_clk_i;
 wire clknet_4_9_0_wb_clk_i;
 wire clknet_4_10_0_wb_clk_i;
 wire clknet_4_11_0_wb_clk_i;
 wire clknet_4_12_0_wb_clk_i;
 wire clknet_4_13_0_wb_clk_i;
 wire clknet_4_14_0_wb_clk_i;
 wire clknet_4_15_0_wb_clk_i;

 sky130_fd_sc_hd__buf_6 _1665_ (.A(net1),
    .X(_1072_));
 sky130_fd_sc_hd__buf_12 _1666_ (.A(_1072_),
    .X(_1073_));
 sky130_fd_sc_hd__clkbuf_16 _1667_ (.A(_1073_),
    .X(_1074_));
 sky130_fd_sc_hd__inv_2 _1668_ (.A(_1074_),
    .Y(_1470_));
 sky130_fd_sc_hd__inv_2 _1669_ (.A(_1074_),
    .Y(_1454_));
 sky130_fd_sc_hd__inv_2 _1670_ (.A(_1074_),
    .Y(_1472_));
 sky130_fd_sc_hd__inv_2 _1671_ (.A(_1074_),
    .Y(_1473_));
 sky130_fd_sc_hd__inv_2 _1672_ (.A(_1074_),
    .Y(_1471_));
 sky130_fd_sc_hd__inv_2 _1673_ (.A(_1074_),
    .Y(_1478_));
 sky130_fd_sc_hd__inv_2 _1674_ (.A(_1074_),
    .Y(_1475_));
 sky130_fd_sc_hd__inv_2 _1675_ (.A(_1074_),
    .Y(_1474_));
 sky130_fd_sc_hd__inv_2 _1676_ (.A(_1074_),
    .Y(_1481_));
 sky130_fd_sc_hd__inv_2 _1677_ (.A(_1074_),
    .Y(_1511_));
 sky130_fd_sc_hd__buf_12 _1678_ (.A(_1073_),
    .X(_1075_));
 sky130_fd_sc_hd__inv_2 _1679_ (.A(_1075_),
    .Y(_1483_));
 sky130_fd_sc_hd__inv_2 _1680_ (.A(_1075_),
    .Y(_1469_));
 sky130_fd_sc_hd__inv_2 _1681_ (.A(_1075_),
    .Y(_1484_));
 sky130_fd_sc_hd__inv_2 _1682_ (.A(_1075_),
    .Y(_1467_));
 sky130_fd_sc_hd__inv_2 _1683_ (.A(_1075_),
    .Y(_1485_));
 sky130_fd_sc_hd__inv_2 _1684_ (.A(_1075_),
    .Y(_1487_));
 sky130_fd_sc_hd__inv_2 _1685_ (.A(_1075_),
    .Y(_1512_));
 sky130_fd_sc_hd__inv_2 _1686_ (.A(_1075_),
    .Y(_1488_));
 sky130_fd_sc_hd__inv_2 _1687_ (.A(_1075_),
    .Y(_1489_));
 sky130_fd_sc_hd__inv_2 _1688_ (.A(_1075_),
    .Y(_1466_));
 sky130_fd_sc_hd__buf_12 _1689_ (.A(_1072_),
    .X(_1076_));
 sky130_fd_sc_hd__inv_2 _1690_ (.A(_1076_),
    .Y(_1455_));
 sky130_fd_sc_hd__inv_2 _1691_ (.A(_1076_),
    .Y(_1463_));
 sky130_fd_sc_hd__inv_2 _1692_ (.A(_1076_),
    .Y(_1476_));
 sky130_fd_sc_hd__inv_2 _1693_ (.A(_1076_),
    .Y(_1477_));
 sky130_fd_sc_hd__inv_2 _1694_ (.A(_1076_),
    .Y(_1465_));
 sky130_fd_sc_hd__inv_2 _1695_ (.A(_1076_),
    .Y(_1464_));
 sky130_fd_sc_hd__inv_2 _1696_ (.A(_1076_),
    .Y(_1490_));
 sky130_fd_sc_hd__inv_2 _1697_ (.A(_1076_),
    .Y(_1491_));
 sky130_fd_sc_hd__inv_2 _1698_ (.A(_1076_),
    .Y(_1492_));
 sky130_fd_sc_hd__inv_2 _1699_ (.A(_1076_),
    .Y(_1459_));
 sky130_fd_sc_hd__clkbuf_16 _1700_ (.A(_1072_),
    .X(_1077_));
 sky130_fd_sc_hd__inv_2 _1701_ (.A(_1077_),
    .Y(_1493_));
 sky130_fd_sc_hd__inv_2 _1702_ (.A(_1077_),
    .Y(_1494_));
 sky130_fd_sc_hd__inv_2 _1703_ (.A(_1077_),
    .Y(_1495_));
 sky130_fd_sc_hd__inv_2 _1704_ (.A(_1077_),
    .Y(_1513_));
 sky130_fd_sc_hd__inv_2 _1705_ (.A(_1077_),
    .Y(_1496_));
 sky130_fd_sc_hd__inv_2 _1706_ (.A(_1077_),
    .Y(_1497_));
 sky130_fd_sc_hd__inv_2 _1707_ (.A(_1077_),
    .Y(_1498_));
 sky130_fd_sc_hd__inv_2 _1708_ (.A(_1077_),
    .Y(_1499_));
 sky130_fd_sc_hd__inv_2 _1709_ (.A(_1077_),
    .Y(_1500_));
 sky130_fd_sc_hd__inv_2 _1710_ (.A(_1077_),
    .Y(_1501_));
 sky130_fd_sc_hd__clkbuf_16 _1711_ (.A(_1072_),
    .X(_1078_));
 sky130_fd_sc_hd__inv_2 _1712_ (.A(_1078_),
    .Y(_1502_));
 sky130_fd_sc_hd__inv_2 _1713_ (.A(_1078_),
    .Y(_1503_));
 sky130_fd_sc_hd__inv_2 _1714_ (.A(_1078_),
    .Y(_1504_));
 sky130_fd_sc_hd__inv_2 _1715_ (.A(_1078_),
    .Y(_1458_));
 sky130_fd_sc_hd__inv_2 _1716_ (.A(_1078_),
    .Y(_1505_));
 sky130_fd_sc_hd__inv_2 _1717_ (.A(_1078_),
    .Y(_1506_));
 sky130_fd_sc_hd__inv_2 _1718_ (.A(_1078_),
    .Y(_1507_));
 sky130_fd_sc_hd__inv_2 _1719_ (.A(_1078_),
    .Y(_1508_));
 sky130_fd_sc_hd__inv_2 _1720_ (.A(_1078_),
    .Y(_1509_));
 sky130_fd_sc_hd__inv_2 _1721_ (.A(_1078_),
    .Y(_1510_));
 sky130_fd_sc_hd__clkbuf_16 _1722_ (.A(_1072_),
    .X(_1079_));
 sky130_fd_sc_hd__inv_2 _1723_ (.A(_1079_),
    .Y(_1482_));
 sky130_fd_sc_hd__inv_2 _1724_ (.A(_1079_),
    .Y(_1515_));
 sky130_fd_sc_hd__inv_2 _1725_ (.A(_1079_),
    .Y(_1516_));
 sky130_fd_sc_hd__inv_2 _1726_ (.A(_1079_),
    .Y(_1517_));
 sky130_fd_sc_hd__inv_2 _1727_ (.A(_1079_),
    .Y(_1518_));
 sky130_fd_sc_hd__inv_2 _1728_ (.A(_1079_),
    .Y(_1519_));
 sky130_fd_sc_hd__inv_2 _1729_ (.A(_1079_),
    .Y(_1520_));
 sky130_fd_sc_hd__inv_2 _1730_ (.A(_1079_),
    .Y(_1521_));
 sky130_fd_sc_hd__inv_2 _1731_ (.A(_1079_),
    .Y(_1522_));
 sky130_fd_sc_hd__inv_2 _1732_ (.A(_1079_),
    .Y(_1523_));
 sky130_fd_sc_hd__buf_12 _1733_ (.A(_1072_),
    .X(_1080_));
 sky130_fd_sc_hd__inv_2 _1734_ (.A(_1080_),
    .Y(_1525_));
 sky130_fd_sc_hd__inv_2 _1735_ (.A(_1080_),
    .Y(_1526_));
 sky130_fd_sc_hd__inv_2 _1736_ (.A(_1080_),
    .Y(_1527_));
 sky130_fd_sc_hd__inv_2 _1737_ (.A(_1080_),
    .Y(_1528_));
 sky130_fd_sc_hd__inv_2 _1738_ (.A(_1080_),
    .Y(_1529_));
 sky130_fd_sc_hd__inv_2 _1739_ (.A(_1080_),
    .Y(_1530_));
 sky130_fd_sc_hd__inv_2 _1740_ (.A(_1080_),
    .Y(_1531_));
 sky130_fd_sc_hd__inv_2 _1741_ (.A(_1080_),
    .Y(_1532_));
 sky130_fd_sc_hd__inv_2 _1742_ (.A(_1080_),
    .Y(_1533_));
 sky130_fd_sc_hd__inv_2 _1743_ (.A(_1080_),
    .Y(_1534_));
 sky130_fd_sc_hd__buf_12 _1744_ (.A(_1072_),
    .X(_1081_));
 sky130_fd_sc_hd__inv_2 _1745_ (.A(_1081_),
    .Y(_1535_));
 sky130_fd_sc_hd__inv_2 _1746_ (.A(_1081_),
    .Y(_1536_));
 sky130_fd_sc_hd__inv_2 _1747_ (.A(_1081_),
    .Y(_1537_));
 sky130_fd_sc_hd__inv_2 _1748_ (.A(_1081_),
    .Y(_1538_));
 sky130_fd_sc_hd__inv_2 _1749_ (.A(_1081_),
    .Y(_1539_));
 sky130_fd_sc_hd__inv_2 _1750_ (.A(_1081_),
    .Y(_1540_));
 sky130_fd_sc_hd__inv_2 _1751_ (.A(_1081_),
    .Y(_1541_));
 sky130_fd_sc_hd__inv_2 _1752_ (.A(_1081_),
    .Y(_1542_));
 sky130_fd_sc_hd__inv_2 _1753_ (.A(_1081_),
    .Y(_1543_));
 sky130_fd_sc_hd__inv_2 _1754_ (.A(_1081_),
    .Y(_1544_));
 sky130_fd_sc_hd__buf_12 _1755_ (.A(_1072_),
    .X(_1082_));
 sky130_fd_sc_hd__inv_2 _1756_ (.A(_1082_),
    .Y(_1545_));
 sky130_fd_sc_hd__inv_2 _1757_ (.A(_1082_),
    .Y(_1546_));
 sky130_fd_sc_hd__inv_2 _1758_ (.A(_1082_),
    .Y(_1547_));
 sky130_fd_sc_hd__inv_2 _1759_ (.A(_1082_),
    .Y(_1548_));
 sky130_fd_sc_hd__inv_2 _1760_ (.A(_1082_),
    .Y(_1549_));
 sky130_fd_sc_hd__inv_2 _1761_ (.A(_1082_),
    .Y(_1550_));
 sky130_fd_sc_hd__inv_2 _1762_ (.A(_1082_),
    .Y(_1551_));
 sky130_fd_sc_hd__inv_2 _1763_ (.A(_1082_),
    .Y(_1552_));
 sky130_fd_sc_hd__inv_2 _1764_ (.A(_1082_),
    .Y(_1553_));
 sky130_fd_sc_hd__inv_2 _1765_ (.A(_1082_),
    .Y(_1554_));
 sky130_fd_sc_hd__buf_8 _1766_ (.A(_1072_),
    .X(_1083_));
 sky130_fd_sc_hd__inv_2 _1767_ (.A(_1083_),
    .Y(_1555_));
 sky130_fd_sc_hd__inv_2 _1768_ (.A(_1083_),
    .Y(_1556_));
 sky130_fd_sc_hd__inv_2 _1769_ (.A(_1083_),
    .Y(_1557_));
 sky130_fd_sc_hd__inv_2 _1770_ (.A(_1083_),
    .Y(_1558_));
 sky130_fd_sc_hd__inv_2 _1771_ (.A(_1083_),
    .Y(_1559_));
 sky130_fd_sc_hd__inv_2 _1772_ (.A(_1083_),
    .Y(_1560_));
 sky130_fd_sc_hd__inv_2 _1773_ (.A(_1083_),
    .Y(_1561_));
 sky130_fd_sc_hd__inv_2 _1774_ (.A(_1083_),
    .Y(_1468_));
 sky130_fd_sc_hd__inv_2 _1775_ (.A(_1083_),
    .Y(_1457_));
 sky130_fd_sc_hd__inv_2 _1776_ (.A(_1083_),
    .Y(_1456_));
 sky130_fd_sc_hd__inv_2 _1777_ (.A(_1073_),
    .Y(_1480_));
 sky130_fd_sc_hd__inv_2 _1778_ (.A(_1073_),
    .Y(_1462_));
 sky130_fd_sc_hd__inv_2 _1779_ (.A(_1073_),
    .Y(_1461_));
 sky130_fd_sc_hd__inv_2 _1780_ (.A(_1073_),
    .Y(_1460_));
 sky130_fd_sc_hd__inv_2 _1781_ (.A(_1073_),
    .Y(_1479_));
 sky130_fd_sc_hd__inv_2 _1782_ (.A(_1073_),
    .Y(_1514_));
 sky130_fd_sc_hd__inv_2 _1783_ (.A(_1073_),
    .Y(_1524_));
 sky130_fd_sc_hd__inv_2 _1784_ (.A(_1073_),
    .Y(_1486_));
 sky130_fd_sc_hd__clkinv_4 _1785_ (.A(net4),
    .Y(_1084_));
 sky130_fd_sc_hd__clkbuf_4 _1786_ (.A(\simon0.state[6] ),
    .X(_1085_));
 sky130_fd_sc_hd__buf_2 _1787_ (.A(\simon0.seq_length[3] ),
    .X(_1086_));
 sky130_fd_sc_hd__and3_1 _1788_ (.A(\simon0.seq_counter[2] ),
    .B(\simon0.seq_counter[1] ),
    .C(\simon0.seq_counter[0] ),
    .X(_1087_));
 sky130_fd_sc_hd__and2_1 _1789_ (.A(\simon0.seq_counter[3] ),
    .B(_1087_),
    .X(_1088_));
 sky130_fd_sc_hd__nor2_1 _1790_ (.A(\simon0.seq_counter[3] ),
    .B(_1087_),
    .Y(_1089_));
 sky130_fd_sc_hd__or2_1 _1791_ (.A(_1088_),
    .B(_1089_),
    .X(_1090_));
 sky130_fd_sc_hd__nand2_1 _1792_ (.A(_1086_),
    .B(_1090_),
    .Y(_1091_));
 sky130_fd_sc_hd__nor2_1 _1793_ (.A(\simon0.seq_counter[4] ),
    .B(_1088_),
    .Y(_1092_));
 sky130_fd_sc_hd__o22a_1 _1794_ (.A1(\simon0.seq_length[3] ),
    .A2(_1090_),
    .B1(_1092_),
    .B2(\simon0.seq_length[4] ),
    .X(_1093_));
 sky130_fd_sc_hd__a21oi_1 _1795_ (.A1(\simon0.seq_counter[1] ),
    .A2(\simon0.seq_counter[0] ),
    .B1(\simon0.seq_counter[2] ),
    .Y(_1094_));
 sky130_fd_sc_hd__or2_1 _1796_ (.A(_1087_),
    .B(_1094_),
    .X(_1095_));
 sky130_fd_sc_hd__nand2_1 _1797_ (.A(\simon0.seq_counter[4] ),
    .B(_1088_),
    .Y(_1096_));
 sky130_fd_sc_hd__a21boi_1 _1798_ (.A1(\simon0.seq_length[2] ),
    .A2(_1095_),
    .B1_N(_1096_),
    .Y(_1097_));
 sky130_fd_sc_hd__xnor2_1 _1799_ (.A(\simon0.seq_counter[1] ),
    .B(\simon0.seq_counter[0] ),
    .Y(_1098_));
 sky130_fd_sc_hd__xnor2_1 _1800_ (.A(\simon0.seq_counter[0] ),
    .B(\simon0.seq_length[0] ),
    .Y(_1099_));
 sky130_fd_sc_hd__a21oi_1 _1801_ (.A1(\simon0.seq_length[1] ),
    .A2(_1098_),
    .B1(_1099_),
    .Y(_1100_));
 sky130_fd_sc_hd__nand2_1 _1802_ (.A(\simon0.seq_length[4] ),
    .B(_1092_),
    .Y(_1101_));
 sky130_fd_sc_hd__o211a_1 _1803_ (.A1(\simon0.seq_length[1] ),
    .A2(_1098_),
    .B1(_1100_),
    .C1(_1101_),
    .X(_1102_));
 sky130_fd_sc_hd__o211a_1 _1804_ (.A1(\simon0.seq_length[2] ),
    .A2(_1095_),
    .B1(_1097_),
    .C1(_1102_),
    .X(_1103_));
 sky130_fd_sc_hd__nand3_4 _1805_ (.A(_1091_),
    .B(_1093_),
    .C(_1103_),
    .Y(_1104_));
 sky130_fd_sc_hd__or4bb_1 _1806_ (.A(\simon0.millis_counter[5] ),
    .B(\simon0.millis_counter[6] ),
    .C_N(\simon0.millis_counter[7] ),
    .D_N(\simon0.millis_counter[4] ),
    .X(_1105_));
 sky130_fd_sc_hd__or2_2 _1807_ (.A(\simon0.millis_counter[0] ),
    .B(\simon0.millis_counter[1] ),
    .X(_1106_));
 sky130_fd_sc_hd__or2_1 _1808_ (.A(\simon0.millis_counter[2] ),
    .B(_1106_),
    .X(_1107_));
 sky130_fd_sc_hd__inv_2 _1809_ (.A(\simon0.millis_counter[9] ),
    .Y(_1108_));
 sky130_fd_sc_hd__nand2_1 _1810_ (.A(\simon0.millis_counter[8] ),
    .B(_1108_),
    .Y(_1109_));
 sky130_fd_sc_hd__or4_2 _1811_ (.A(\simon0.millis_counter[3] ),
    .B(_1105_),
    .C(_1107_),
    .D(_1109_),
    .X(_1110_));
 sky130_fd_sc_hd__inv_2 _1812_ (.A(_1110_),
    .Y(_1111_));
 sky130_fd_sc_hd__buf_2 _1813_ (.A(\simon0.state[3] ),
    .X(_1112_));
 sky130_fd_sc_hd__or3b_1 _1814_ (.A(\simon0.millis_counter[0] ),
    .B(\simon0.millis_counter[3] ),
    .C_N(\simon0.millis_counter[2] ),
    .X(_1113_));
 sky130_fd_sc_hd__or4b_1 _1815_ (.A(\simon0.millis_counter[8] ),
    .B(\simon0.millis_counter[9] ),
    .C(_1105_),
    .D_N(\simon0.millis_counter[1] ),
    .X(_1114_));
 sky130_fd_sc_hd__nor2_1 _1816_ (.A(_1113_),
    .B(_1114_),
    .Y(_1115_));
 sky130_fd_sc_hd__and3_1 _1817_ (.A(\simon0.tone_sequence_counter[0] ),
    .B(\simon0.tone_sequence_counter[1] ),
    .C(\simon0.tone_sequence_counter[2] ),
    .X(_1116_));
 sky130_fd_sc_hd__and4_1 _1818_ (.A(\simon0.millis_counter[4] ),
    .B(\simon0.millis_counter[5] ),
    .C(\simon0.millis_counter[6] ),
    .D(\simon0.millis_counter[7] ),
    .X(_1117_));
 sky130_fd_sc_hd__or3b_1 _1819_ (.A(\simon0.millis_counter[1] ),
    .B(_1109_),
    .C_N(_1117_),
    .X(_1118_));
 sky130_fd_sc_hd__nor2_1 _1820_ (.A(_1113_),
    .B(_1118_),
    .Y(_1119_));
 sky130_fd_sc_hd__a32o_1 _1821_ (.A1(_1112_),
    .A2(_1115_),
    .A3(_1116_),
    .B1(_1119_),
    .B2(\simon0.state[4] ),
    .X(_1120_));
 sky130_fd_sc_hd__a31o_1 _1822_ (.A1(_1085_),
    .A2(_1104_),
    .A3(_1111_),
    .B1(_1120_),
    .X(_1121_));
 sky130_fd_sc_hd__and2_1 _1823_ (.A(_1084_),
    .B(_1121_),
    .X(_1122_));
 sky130_fd_sc_hd__clkbuf_1 _1824_ (.A(_1122_),
    .X(_0007_));
 sky130_fd_sc_hd__clkbuf_4 _1825_ (.A(net4),
    .X(_1123_));
 sky130_fd_sc_hd__clkbuf_4 _1826_ (.A(_1123_),
    .X(_1124_));
 sky130_fd_sc_hd__inv_2 _1827_ (.A(\simon0.user_input[0] ),
    .Y(_1125_));
 sky130_fd_sc_hd__inv_2 _1828_ (.A(_0003_),
    .Y(_1126_));
 sky130_fd_sc_hd__mux4_1 _1829_ (.A0(\simon0.seq[20][0] ),
    .A1(\simon0.seq[21][0] ),
    .A2(\simon0.seq[22][0] ),
    .A3(\simon0.seq[23][0] ),
    .S0(_0000_),
    .S1(_0001_),
    .X(_1127_));
 sky130_fd_sc_hd__mux4_1 _1830_ (.A0(\simon0.seq[16][0] ),
    .A1(\simon0.seq[17][0] ),
    .A2(\simon0.seq[18][0] ),
    .A3(\simon0.seq[19][0] ),
    .S0(_0000_),
    .S1(_0001_),
    .X(_1128_));
 sky130_fd_sc_hd__clkinv_2 _1831_ (.A(_0002_),
    .Y(_1129_));
 sky130_fd_sc_hd__mux2_1 _1832_ (.A0(_1127_),
    .A1(_1128_),
    .S(_1129_),
    .X(_1130_));
 sky130_fd_sc_hd__buf_4 _1833_ (.A(_0000_),
    .X(_1131_));
 sky130_fd_sc_hd__clkbuf_4 _1834_ (.A(_0001_),
    .X(_1132_));
 sky130_fd_sc_hd__mux4_1 _1835_ (.A0(\simon0.seq[24][0] ),
    .A1(\simon0.seq[25][0] ),
    .A2(\simon0.seq[26][0] ),
    .A3(\simon0.seq[27][0] ),
    .S0(_1131_),
    .S1(_1132_),
    .X(_1133_));
 sky130_fd_sc_hd__or2_1 _1836_ (.A(_0002_),
    .B(_1133_),
    .X(_1134_));
 sky130_fd_sc_hd__mux4_1 _1837_ (.A0(\simon0.seq[28][0] ),
    .A1(\simon0.seq[29][0] ),
    .A2(\simon0.seq[30][0] ),
    .A3(\simon0.seq[31][0] ),
    .S0(_1131_),
    .S1(_1132_),
    .X(_1135_));
 sky130_fd_sc_hd__o21a_1 _1838_ (.A1(_1129_),
    .A2(_1135_),
    .B1(_0003_),
    .X(_1136_));
 sky130_fd_sc_hd__inv_2 _1839_ (.A(_0004_),
    .Y(_1137_));
 sky130_fd_sc_hd__a221o_1 _1840_ (.A1(_1126_),
    .A2(_1130_),
    .B1(_1134_),
    .B2(_1136_),
    .C1(_1137_),
    .X(_1138_));
 sky130_fd_sc_hd__mux4_1 _1841_ (.A0(\simon0.seq[8][0] ),
    .A1(\simon0.seq[9][0] ),
    .A2(\simon0.seq[10][0] ),
    .A3(\simon0.seq[11][0] ),
    .S0(_1131_),
    .S1(_1132_),
    .X(_1139_));
 sky130_fd_sc_hd__or2_1 _1842_ (.A(_0002_),
    .B(_1139_),
    .X(_1140_));
 sky130_fd_sc_hd__mux4_1 _1843_ (.A0(\simon0.seq[12][0] ),
    .A1(\simon0.seq[13][0] ),
    .A2(\simon0.seq[14][0] ),
    .A3(\simon0.seq[15][0] ),
    .S0(_1131_),
    .S1(_1132_),
    .X(_1141_));
 sky130_fd_sc_hd__o21a_1 _1844_ (.A1(_1129_),
    .A2(_1141_),
    .B1(_0003_),
    .X(_1142_));
 sky130_fd_sc_hd__mux4_1 _1845_ (.A0(\simon0.seq[4][0] ),
    .A1(\simon0.seq[5][0] ),
    .A2(\simon0.seq[6][0] ),
    .A3(\simon0.seq[7][0] ),
    .S0(_1131_),
    .S1(_1132_),
    .X(_1143_));
 sky130_fd_sc_hd__mux4_1 _1846_ (.A0(\simon0.seq[0][0] ),
    .A1(\simon0.seq[1][0] ),
    .A2(\simon0.seq[2][0] ),
    .A3(\simon0.seq[3][0] ),
    .S0(_1131_),
    .S1(_1132_),
    .X(_1144_));
 sky130_fd_sc_hd__mux2_1 _1847_ (.A0(_1143_),
    .A1(_1144_),
    .S(_1129_),
    .X(_1145_));
 sky130_fd_sc_hd__a221o_1 _1848_ (.A1(_1140_),
    .A2(_1142_),
    .B1(_1145_),
    .B2(_1126_),
    .C1(_0004_),
    .X(_1146_));
 sky130_fd_sc_hd__nand2_1 _1849_ (.A(_1138_),
    .B(_1146_),
    .Y(_1147_));
 sky130_fd_sc_hd__xnor2_1 _1850_ (.A(_1125_),
    .B(_1147_),
    .Y(_1148_));
 sky130_fd_sc_hd__inv_2 _1851_ (.A(\simon0.user_input[1] ),
    .Y(_1149_));
 sky130_fd_sc_hd__mux4_1 _1852_ (.A0(\simon0.seq[20][1] ),
    .A1(\simon0.seq[21][1] ),
    .A2(\simon0.seq[22][1] ),
    .A3(\simon0.seq[23][1] ),
    .S0(_0000_),
    .S1(_0001_),
    .X(_1150_));
 sky130_fd_sc_hd__mux4_1 _1853_ (.A0(\simon0.seq[16][1] ),
    .A1(\simon0.seq[17][1] ),
    .A2(\simon0.seq[18][1] ),
    .A3(\simon0.seq[19][1] ),
    .S0(_0000_),
    .S1(_0001_),
    .X(_1151_));
 sky130_fd_sc_hd__mux2_1 _1854_ (.A0(_1150_),
    .A1(_1151_),
    .S(_1129_),
    .X(_1152_));
 sky130_fd_sc_hd__mux4_1 _1855_ (.A0(\simon0.seq[24][1] ),
    .A1(\simon0.seq[25][1] ),
    .A2(\simon0.seq[26][1] ),
    .A3(\simon0.seq[27][1] ),
    .S0(_1131_),
    .S1(_1132_),
    .X(_1153_));
 sky130_fd_sc_hd__or2_1 _1856_ (.A(_0002_),
    .B(_1153_),
    .X(_1154_));
 sky130_fd_sc_hd__mux4_1 _1857_ (.A0(\simon0.seq[28][1] ),
    .A1(\simon0.seq[29][1] ),
    .A2(\simon0.seq[30][1] ),
    .A3(\simon0.seq[31][1] ),
    .S0(_1131_),
    .S1(_1132_),
    .X(_1155_));
 sky130_fd_sc_hd__o21a_1 _1858_ (.A1(_1129_),
    .A2(_1155_),
    .B1(_0003_),
    .X(_1156_));
 sky130_fd_sc_hd__a221o_1 _1859_ (.A1(_1126_),
    .A2(_1152_),
    .B1(_1154_),
    .B2(_1156_),
    .C1(_1137_),
    .X(_1157_));
 sky130_fd_sc_hd__mux4_1 _1860_ (.A0(\simon0.seq[4][1] ),
    .A1(\simon0.seq[5][1] ),
    .A2(\simon0.seq[6][1] ),
    .A3(\simon0.seq[7][1] ),
    .S0(_0000_),
    .S1(_0001_),
    .X(_1158_));
 sky130_fd_sc_hd__mux4_1 _1861_ (.A0(\simon0.seq[0][1] ),
    .A1(\simon0.seq[1][1] ),
    .A2(\simon0.seq[2][1] ),
    .A3(\simon0.seq[3][1] ),
    .S0(_0000_),
    .S1(_0001_),
    .X(_1159_));
 sky130_fd_sc_hd__mux2_1 _1862_ (.A0(_1158_),
    .A1(_1159_),
    .S(_1129_),
    .X(_1160_));
 sky130_fd_sc_hd__mux4_1 _1863_ (.A0(\simon0.seq[8][1] ),
    .A1(\simon0.seq[9][1] ),
    .A2(\simon0.seq[10][1] ),
    .A3(\simon0.seq[11][1] ),
    .S0(_1131_),
    .S1(_1132_),
    .X(_1161_));
 sky130_fd_sc_hd__or2_1 _1864_ (.A(_0002_),
    .B(_1161_),
    .X(_1162_));
 sky130_fd_sc_hd__mux4_1 _1865_ (.A0(\simon0.seq[12][1] ),
    .A1(\simon0.seq[13][1] ),
    .A2(\simon0.seq[14][1] ),
    .A3(\simon0.seq[15][1] ),
    .S0(_1131_),
    .S1(_1132_),
    .X(_1163_));
 sky130_fd_sc_hd__o21a_1 _1866_ (.A1(_1129_),
    .A2(_1163_),
    .B1(_0003_),
    .X(_1164_));
 sky130_fd_sc_hd__a221o_1 _1867_ (.A1(_1126_),
    .A2(_1160_),
    .B1(_1162_),
    .B2(_1164_),
    .C1(_0004_),
    .X(_1165_));
 sky130_fd_sc_hd__nand2_1 _1868_ (.A(_1157_),
    .B(_1165_),
    .Y(_1166_));
 sky130_fd_sc_hd__xnor2_1 _1869_ (.A(_1149_),
    .B(_1166_),
    .Y(_1167_));
 sky130_fd_sc_hd__and3_1 _1870_ (.A(_1104_),
    .B(_1148_),
    .C(_1167_),
    .X(_1168_));
 sky130_fd_sc_hd__buf_4 _1871_ (.A(\simon0.state[5] ),
    .X(_1169_));
 sky130_fd_sc_hd__inv_2 _1872_ (.A(_1169_),
    .Y(_1170_));
 sky130_fd_sc_hd__or4bb_1 _1873_ (.A(\simon0.millis_counter[6] ),
    .B(\simon0.millis_counter[7] ),
    .C_N(\simon0.millis_counter[2] ),
    .D_N(\simon0.millis_counter[3] ),
    .X(_1171_));
 sky130_fd_sc_hd__or2b_1 _1874_ (.A(\simon0.millis_counter[4] ),
    .B_N(\simon0.millis_counter[5] ),
    .X(_1172_));
 sky130_fd_sc_hd__or4_4 _1875_ (.A(_1106_),
    .B(_1109_),
    .C(_1171_),
    .D(_1172_),
    .X(_1173_));
 sky130_fd_sc_hd__nor2_1 _1876_ (.A(_1170_),
    .B(_1173_),
    .Y(_1174_));
 sky130_fd_sc_hd__or2_1 _1877_ (.A(net6),
    .B(net2),
    .X(_1175_));
 sky130_fd_sc_hd__a21oi_1 _1878_ (.A1(net7),
    .A2(net3),
    .B1(_1175_),
    .Y(_1176_));
 sky130_fd_sc_hd__o21a_1 _1879_ (.A1(net7),
    .A2(net3),
    .B1(_1176_),
    .X(_1177_));
 sky130_fd_sc_hd__or3b_1 _1880_ (.A(net7),
    .B(net3),
    .C_N(_1175_),
    .X(_1178_));
 sky130_fd_sc_hd__a21oi_1 _1881_ (.A1(net6),
    .A2(net2),
    .B1(_1178_),
    .Y(_1179_));
 sky130_fd_sc_hd__nor2_1 _1882_ (.A(_1177_),
    .B(_1179_),
    .Y(_1180_));
 sky130_fd_sc_hd__nor2_1 _1883_ (.A(_1104_),
    .B(_1110_),
    .Y(_1181_));
 sky130_fd_sc_hd__a22o_1 _1884_ (.A1(\simon0.state[1] ),
    .A2(_1180_),
    .B1(_1181_),
    .B2(_1085_),
    .X(_1182_));
 sky130_fd_sc_hd__a21oi_1 _1885_ (.A1(_1168_),
    .A2(_1174_),
    .B1(_1182_),
    .Y(_1183_));
 sky130_fd_sc_hd__nor2_1 _1886_ (.A(_1124_),
    .B(_1183_),
    .Y(_0006_));
 sky130_fd_sc_hd__nor3_4 _1887_ (.A(net7),
    .B(net3),
    .C(_1175_),
    .Y(_1184_));
 sky130_fd_sc_hd__a21o_1 _1888_ (.A1(\simon0.state[0] ),
    .A2(_1184_),
    .B1(_1124_),
    .X(_0005_));
 sky130_fd_sc_hd__nand2_1 _1889_ (.A(_1148_),
    .B(_1167_),
    .Y(_1185_));
 sky130_fd_sc_hd__and2_1 _1890_ (.A(\simon0.state[7] ),
    .B(_1184_),
    .X(_1186_));
 sky130_fd_sc_hd__buf_2 _1891_ (.A(_1186_),
    .X(_1187_));
 sky130_fd_sc_hd__a21oi_1 _1892_ (.A1(_1185_),
    .A2(_1174_),
    .B1(_1187_),
    .Y(_1188_));
 sky130_fd_sc_hd__nor2_1 _1893_ (.A(_1124_),
    .B(_1188_),
    .Y(_0012_));
 sky130_fd_sc_hd__and2_1 _1894_ (.A(_1085_),
    .B(_1110_),
    .X(_1189_));
 sky130_fd_sc_hd__clkbuf_4 _1895_ (.A(_1084_),
    .X(_1190_));
 sky130_fd_sc_hd__o21a_1 _1896_ (.A1(\simon0.state[2] ),
    .A2(_1189_),
    .B1(_1190_),
    .X(_0011_));
 sky130_fd_sc_hd__and2_1 _1897_ (.A(_1169_),
    .B(_1173_),
    .X(_1191_));
 sky130_fd_sc_hd__nor2_1 _1898_ (.A(net4),
    .B(_1184_),
    .Y(_1192_));
 sky130_fd_sc_hd__o211a_1 _1899_ (.A1(_1177_),
    .A2(_1179_),
    .B1(_1192_),
    .C1(\simon0.state[1] ),
    .X(_1193_));
 sky130_fd_sc_hd__a21o_1 _1900_ (.A1(_1190_),
    .A2(_1191_),
    .B1(_1193_),
    .X(_0010_));
 sky130_fd_sc_hd__clkbuf_4 _1901_ (.A(_1084_),
    .X(_1194_));
 sky130_fd_sc_hd__or2_1 _1902_ (.A(_1113_),
    .B(_1118_),
    .X(_1195_));
 sky130_fd_sc_hd__or2_1 _1903_ (.A(\simon0.state[0] ),
    .B(\simon0.state[7] ),
    .X(_1196_));
 sky130_fd_sc_hd__a32o_1 _1904_ (.A1(\simon0.state[4] ),
    .A2(_1194_),
    .A3(_1195_),
    .B1(_1192_),
    .B2(_1196_),
    .X(_0009_));
 sky130_fd_sc_hd__inv_2 _1905_ (.A(_1112_),
    .Y(_1197_));
 sky130_fd_sc_hd__a21o_1 _1906_ (.A1(_1115_),
    .A2(_1116_),
    .B1(_1197_),
    .X(_1198_));
 sky130_fd_sc_hd__or3_1 _1907_ (.A(_1170_),
    .B(_1185_),
    .C(_1173_),
    .X(_1199_));
 sky130_fd_sc_hd__or2_1 _1908_ (.A(_1104_),
    .B(_1199_),
    .X(_1200_));
 sky130_fd_sc_hd__buf_4 _1909_ (.A(_1123_),
    .X(_1201_));
 sky130_fd_sc_hd__a21oi_1 _1910_ (.A1(_1198_),
    .A2(_1200_),
    .B1(_1201_),
    .Y(_0008_));
 sky130_fd_sc_hd__or4_1 _1911_ (.A(\simon0.state[3] ),
    .B(\simon0.state[1] ),
    .C(\simon0.state[0] ),
    .D(\simon0.state[2] ),
    .X(_1202_));
 sky130_fd_sc_hd__or3_1 _1912_ (.A(\simon0.state[6] ),
    .B(\simon0.state[3] ),
    .C(\simon0.state[5] ),
    .X(_1203_));
 sky130_fd_sc_hd__or2_1 _1913_ (.A(\simon0.state[7] ),
    .B(_1203_),
    .X(_1204_));
 sky130_fd_sc_hd__buf_2 _1914_ (.A(_1204_),
    .X(_1205_));
 sky130_fd_sc_hd__nor2_1 _1915_ (.A(_1202_),
    .B(_1205_),
    .Y(_1206_));
 sky130_fd_sc_hd__or4_1 _1916_ (.A(\simon0.state[4] ),
    .B(net4),
    .C(\simon0.state[6] ),
    .D(\simon0.state[7] ),
    .X(_1207_));
 sky130_fd_sc_hd__or4_1 _1917_ (.A(_1104_),
    .B(_1173_),
    .C(_1202_),
    .D(_1207_),
    .X(_1208_));
 sky130_fd_sc_hd__nor2_1 _1918_ (.A(_1185_),
    .B(_1208_),
    .Y(_1209_));
 sky130_fd_sc_hd__buf_2 _1919_ (.A(_1209_),
    .X(_1210_));
 sky130_fd_sc_hd__a21o_1 _1920_ (.A1(_1084_),
    .A2(_1206_),
    .B1(_1210_),
    .X(_1211_));
 sky130_fd_sc_hd__and2_2 _1921_ (.A(\simon0.next_random[0] ),
    .B(_1211_),
    .X(_1212_));
 sky130_fd_sc_hd__buf_2 _1922_ (.A(_1212_),
    .X(_1213_));
 sky130_fd_sc_hd__nand2_1 _1923_ (.A(\simon0.seq_length[0] ),
    .B(_1209_),
    .Y(_1214_));
 sky130_fd_sc_hd__nand2_1 _1924_ (.A(\simon0.seq_length[1] ),
    .B(_1209_),
    .Y(_1215_));
 sky130_fd_sc_hd__and2_1 _1925_ (.A(_1214_),
    .B(_1215_),
    .X(_1216_));
 sky130_fd_sc_hd__buf_2 _1926_ (.A(\simon0.seq_length[4] ),
    .X(_1217_));
 sky130_fd_sc_hd__buf_2 _1927_ (.A(\simon0.seq_length[2] ),
    .X(_1218_));
 sky130_fd_sc_hd__and4b_1 _1928_ (.A_N(_1217_),
    .B(_1086_),
    .C(_1218_),
    .D(_1210_),
    .X(_1219_));
 sky130_fd_sc_hd__nand2_1 _1929_ (.A(_1216_),
    .B(_1219_),
    .Y(_1220_));
 sky130_fd_sc_hd__mux2_1 _1930_ (.A0(_1213_),
    .A1(\simon0.seq[12][0] ),
    .S(_1220_),
    .X(_1221_));
 sky130_fd_sc_hd__clkbuf_1 _1931_ (.A(_1221_),
    .X(_0013_));
 sky130_fd_sc_hd__and2_2 _1932_ (.A(\simon0.next_random[1] ),
    .B(_1211_),
    .X(_1222_));
 sky130_fd_sc_hd__buf_2 _1933_ (.A(_1222_),
    .X(_1223_));
 sky130_fd_sc_hd__mux2_1 _1934_ (.A0(_1223_),
    .A1(\simon0.seq[12][1] ),
    .S(_1220_),
    .X(_1224_));
 sky130_fd_sc_hd__clkbuf_1 _1935_ (.A(_1224_),
    .X(_0014_));
 sky130_fd_sc_hd__nand2_1 _1936_ (.A(_1086_),
    .B(_1210_),
    .Y(_1225_));
 sky130_fd_sc_hd__or3_1 _1937_ (.A(_1217_),
    .B(_1218_),
    .C(_1225_),
    .X(_1226_));
 sky130_fd_sc_hd__nand3_1 _1938_ (.A(\simon0.seq_length[1] ),
    .B(\simon0.seq_length[0] ),
    .C(_1210_),
    .Y(_1227_));
 sky130_fd_sc_hd__or2_1 _1939_ (.A(_1226_),
    .B(_1227_),
    .X(_1228_));
 sky130_fd_sc_hd__mux2_1 _1940_ (.A0(_1213_),
    .A1(\simon0.seq[11][0] ),
    .S(_1228_),
    .X(_1229_));
 sky130_fd_sc_hd__clkbuf_1 _1941_ (.A(_1229_),
    .X(_0015_));
 sky130_fd_sc_hd__mux2_1 _1942_ (.A0(_1223_),
    .A1(\simon0.seq[11][1] ),
    .S(_1228_),
    .X(_1230_));
 sky130_fd_sc_hd__clkbuf_1 _1943_ (.A(_1230_),
    .X(_0016_));
 sky130_fd_sc_hd__buf_2 _1944_ (.A(_1212_),
    .X(_1231_));
 sky130_fd_sc_hd__or2_1 _1945_ (.A(\simon0.seq_length[0] ),
    .B(_1215_),
    .X(_1232_));
 sky130_fd_sc_hd__clkbuf_2 _1946_ (.A(_1232_),
    .X(_1233_));
 sky130_fd_sc_hd__nor2_1 _1947_ (.A(_1226_),
    .B(_1233_),
    .Y(_1234_));
 sky130_fd_sc_hd__mux2_1 _1948_ (.A0(\simon0.seq[10][0] ),
    .A1(_1231_),
    .S(_1234_),
    .X(_1235_));
 sky130_fd_sc_hd__clkbuf_1 _1949_ (.A(_1235_),
    .X(_0017_));
 sky130_fd_sc_hd__buf_2 _1950_ (.A(_1222_),
    .X(_1236_));
 sky130_fd_sc_hd__mux2_1 _1951_ (.A0(\simon0.seq[10][1] ),
    .A1(_1236_),
    .S(_1234_),
    .X(_1237_));
 sky130_fd_sc_hd__clkbuf_1 _1952_ (.A(_1237_),
    .X(_0018_));
 sky130_fd_sc_hd__nand2_2 _1953_ (.A(_1214_),
    .B(_1215_),
    .Y(_1238_));
 sky130_fd_sc_hd__or4bb_2 _1954_ (.A(_1086_),
    .B(\simon0.seq_length[2] ),
    .C_N(_1210_),
    .D_N(_1217_),
    .X(_1239_));
 sky130_fd_sc_hd__nor2_1 _1955_ (.A(_1238_),
    .B(_1239_),
    .Y(_1240_));
 sky130_fd_sc_hd__mux2_1 _1956_ (.A0(\simon0.seq[16][0] ),
    .A1(_1231_),
    .S(_1240_),
    .X(_1241_));
 sky130_fd_sc_hd__clkbuf_1 _1957_ (.A(_1241_),
    .X(_0019_));
 sky130_fd_sc_hd__mux2_1 _1958_ (.A0(\simon0.seq[16][1] ),
    .A1(_1236_),
    .S(_1240_),
    .X(_1242_));
 sky130_fd_sc_hd__clkbuf_1 _1959_ (.A(_1242_),
    .X(_0020_));
 sky130_fd_sc_hd__nor2_1 _1960_ (.A(\simon0.seq_length[1] ),
    .B(_1214_),
    .Y(_1243_));
 sky130_fd_sc_hd__and4_1 _1961_ (.A(_1217_),
    .B(_1086_),
    .C(_1218_),
    .D(_1210_),
    .X(_1244_));
 sky130_fd_sc_hd__nand2_1 _1962_ (.A(_1243_),
    .B(_1244_),
    .Y(_1245_));
 sky130_fd_sc_hd__mux2_1 _1963_ (.A0(_1213_),
    .A1(\simon0.seq[29][0] ),
    .S(_1245_),
    .X(_1246_));
 sky130_fd_sc_hd__clkbuf_1 _1964_ (.A(_1246_),
    .X(_0021_));
 sky130_fd_sc_hd__mux2_1 _1965_ (.A0(_1223_),
    .A1(\simon0.seq[29][1] ),
    .S(_1245_),
    .X(_1247_));
 sky130_fd_sc_hd__clkbuf_1 _1966_ (.A(_1247_),
    .X(_0022_));
 sky130_fd_sc_hd__and3_1 _1967_ (.A(\simon0.seq_length[1] ),
    .B(\simon0.seq_length[0] ),
    .C(_1210_),
    .X(_1248_));
 sky130_fd_sc_hd__nand2_1 _1968_ (.A(_1219_),
    .B(_1248_),
    .Y(_1249_));
 sky130_fd_sc_hd__mux2_1 _1969_ (.A0(_1213_),
    .A1(\simon0.seq[15][0] ),
    .S(_1249_),
    .X(_1250_));
 sky130_fd_sc_hd__clkbuf_1 _1970_ (.A(_1250_),
    .X(_0023_));
 sky130_fd_sc_hd__mux2_1 _1971_ (.A0(_1223_),
    .A1(\simon0.seq[15][1] ),
    .S(_1249_),
    .X(_1251_));
 sky130_fd_sc_hd__clkbuf_1 _1972_ (.A(_1251_),
    .X(_0024_));
 sky130_fd_sc_hd__nor2_1 _1973_ (.A(\simon0.seq_length[0] ),
    .B(_1215_),
    .Y(_1252_));
 sky130_fd_sc_hd__nand2_1 _1974_ (.A(_1219_),
    .B(_1252_),
    .Y(_1253_));
 sky130_fd_sc_hd__mux2_1 _1975_ (.A0(_1213_),
    .A1(\simon0.seq[14][0] ),
    .S(_1253_),
    .X(_1254_));
 sky130_fd_sc_hd__clkbuf_1 _1976_ (.A(_1254_),
    .X(_0025_));
 sky130_fd_sc_hd__mux2_1 _1977_ (.A0(_1223_),
    .A1(\simon0.seq[14][1] ),
    .S(_1253_),
    .X(_1255_));
 sky130_fd_sc_hd__clkbuf_1 _1978_ (.A(_1255_),
    .X(_0026_));
 sky130_fd_sc_hd__nand2_1 _1979_ (.A(_1219_),
    .B(_1243_),
    .Y(_1256_));
 sky130_fd_sc_hd__mux2_1 _1980_ (.A0(_1213_),
    .A1(\simon0.seq[13][0] ),
    .S(_1256_),
    .X(_1257_));
 sky130_fd_sc_hd__clkbuf_1 _1981_ (.A(_1257_),
    .X(_0027_));
 sky130_fd_sc_hd__mux2_1 _1982_ (.A0(_1223_),
    .A1(\simon0.seq[13][1] ),
    .S(_1256_),
    .X(_1258_));
 sky130_fd_sc_hd__clkbuf_1 _1983_ (.A(_1258_),
    .X(_0028_));
 sky130_fd_sc_hd__nor2_1 _1984_ (.A(_1238_),
    .B(_1226_),
    .Y(_1259_));
 sky130_fd_sc_hd__mux2_1 _1985_ (.A0(\simon0.seq[8][0] ),
    .A1(_1231_),
    .S(_1259_),
    .X(_1260_));
 sky130_fd_sc_hd__clkbuf_1 _1986_ (.A(_1260_),
    .X(_0029_));
 sky130_fd_sc_hd__mux2_1 _1987_ (.A0(\simon0.seq[8][1] ),
    .A1(_1236_),
    .S(_1259_),
    .X(_1261_));
 sky130_fd_sc_hd__clkbuf_1 _1988_ (.A(_1261_),
    .X(_0030_));
 sky130_fd_sc_hd__mux2_1 _1989_ (.A0(\simon0.user_input[0] ),
    .A1(_1177_),
    .S(_1193_),
    .X(_1262_));
 sky130_fd_sc_hd__clkbuf_1 _1990_ (.A(_1262_),
    .X(_0031_));
 sky130_fd_sc_hd__nor2_1 _1991_ (.A(net6),
    .B(net7),
    .Y(_1263_));
 sky130_fd_sc_hd__mux2_1 _1992_ (.A0(\simon0.user_input[1] ),
    .A1(_1263_),
    .S(_1193_),
    .X(_1264_));
 sky130_fd_sc_hd__clkbuf_1 _1993_ (.A(_1264_),
    .X(_0032_));
 sky130_fd_sc_hd__nand2_1 _1994_ (.A(\simon0.seq_length[1] ),
    .B(\simon0.seq_length[0] ),
    .Y(_1265_));
 sky130_fd_sc_hd__or4bb_2 _1995_ (.A(_1217_),
    .B(_1086_),
    .C_N(_1218_),
    .D_N(_1210_),
    .X(_1266_));
 sky130_fd_sc_hd__nor2_1 _1996_ (.A(_1265_),
    .B(_1266_),
    .Y(_1267_));
 sky130_fd_sc_hd__mux2_1 _1997_ (.A0(\simon0.seq[7][0] ),
    .A1(_1231_),
    .S(_1267_),
    .X(_1268_));
 sky130_fd_sc_hd__clkbuf_1 _1998_ (.A(_1268_),
    .X(_0033_));
 sky130_fd_sc_hd__mux2_1 _1999_ (.A0(\simon0.seq[7][1] ),
    .A1(_1236_),
    .S(_1267_),
    .X(_1269_));
 sky130_fd_sc_hd__clkbuf_1 _2000_ (.A(_1269_),
    .X(_0034_));
 sky130_fd_sc_hd__nor2_1 _2001_ (.A(_1233_),
    .B(_1266_),
    .Y(_1270_));
 sky130_fd_sc_hd__mux2_1 _2002_ (.A0(\simon0.seq[6][0] ),
    .A1(_1231_),
    .S(_1270_),
    .X(_1271_));
 sky130_fd_sc_hd__clkbuf_1 _2003_ (.A(_1271_),
    .X(_0035_));
 sky130_fd_sc_hd__mux2_1 _2004_ (.A0(\simon0.seq[6][1] ),
    .A1(_1236_),
    .S(_1270_),
    .X(_1272_));
 sky130_fd_sc_hd__clkbuf_1 _2005_ (.A(_1272_),
    .X(_0036_));
 sky130_fd_sc_hd__buf_2 _2006_ (.A(_1212_),
    .X(_1273_));
 sky130_fd_sc_hd__o22a_1 _2007_ (.A1(net4),
    .A2(_1206_),
    .B1(_1208_),
    .B2(_1185_),
    .X(_1274_));
 sky130_fd_sc_hd__mux2_1 _2008_ (.A0(\simon0.seq[0][0] ),
    .A1(_1273_),
    .S(_1274_),
    .X(_1275_));
 sky130_fd_sc_hd__clkbuf_1 _2009_ (.A(_1275_),
    .X(_0037_));
 sky130_fd_sc_hd__buf_2 _2010_ (.A(_1222_),
    .X(_1276_));
 sky130_fd_sc_hd__mux2_1 _2011_ (.A0(\simon0.seq[0][1] ),
    .A1(_1276_),
    .S(_1274_),
    .X(_1277_));
 sky130_fd_sc_hd__clkbuf_1 _2012_ (.A(_1277_),
    .X(_0038_));
 sky130_fd_sc_hd__or2_2 _2013_ (.A(\simon0.seq_length[1] ),
    .B(_1214_),
    .X(_1278_));
 sky130_fd_sc_hd__nor2_1 _2014_ (.A(_1278_),
    .B(_1266_),
    .Y(_1279_));
 sky130_fd_sc_hd__mux2_1 _2015_ (.A0(\simon0.seq[5][0] ),
    .A1(_1273_),
    .S(_1279_),
    .X(_1280_));
 sky130_fd_sc_hd__clkbuf_1 _2016_ (.A(_1280_),
    .X(_0039_));
 sky130_fd_sc_hd__mux2_1 _2017_ (.A0(\simon0.seq[5][1] ),
    .A1(_1276_),
    .S(_1279_),
    .X(_1281_));
 sky130_fd_sc_hd__clkbuf_1 _2018_ (.A(_1281_),
    .X(_0040_));
 sky130_fd_sc_hd__nor2_1 _2019_ (.A(_1238_),
    .B(_1266_),
    .Y(_1282_));
 sky130_fd_sc_hd__mux2_1 _2020_ (.A0(\simon0.seq[4][0] ),
    .A1(_1273_),
    .S(_1282_),
    .X(_1283_));
 sky130_fd_sc_hd__clkbuf_1 _2021_ (.A(_1283_),
    .X(_0041_));
 sky130_fd_sc_hd__mux2_1 _2022_ (.A0(\simon0.seq[4][1] ),
    .A1(_1276_),
    .S(_1282_),
    .X(_1284_));
 sky130_fd_sc_hd__clkbuf_1 _2023_ (.A(_1284_),
    .X(_0042_));
 sky130_fd_sc_hd__o31a_1 _2024_ (.A1(_1217_),
    .A2(_1086_),
    .A3(_1218_),
    .B1(_1210_),
    .X(_1285_));
 sky130_fd_sc_hd__nor2_1 _2025_ (.A(_1227_),
    .B(_1285_),
    .Y(_1286_));
 sky130_fd_sc_hd__mux2_1 _2026_ (.A0(\simon0.seq[3][0] ),
    .A1(_1273_),
    .S(_1286_),
    .X(_1287_));
 sky130_fd_sc_hd__clkbuf_1 _2027_ (.A(_1287_),
    .X(_0043_));
 sky130_fd_sc_hd__mux2_1 _2028_ (.A0(\simon0.seq[3][1] ),
    .A1(_1276_),
    .S(_1286_),
    .X(_1288_));
 sky130_fd_sc_hd__clkbuf_1 _2029_ (.A(_1288_),
    .X(_0044_));
 sky130_fd_sc_hd__and4b_1 _2030_ (.A_N(_1086_),
    .B(_1218_),
    .C(_1210_),
    .D(_1217_),
    .X(_1289_));
 sky130_fd_sc_hd__nand2_1 _2031_ (.A(_1252_),
    .B(_1289_),
    .Y(_1290_));
 sky130_fd_sc_hd__mux2_1 _2032_ (.A0(_1213_),
    .A1(\simon0.seq[22][0] ),
    .S(_1290_),
    .X(_1291_));
 sky130_fd_sc_hd__clkbuf_1 _2033_ (.A(_1291_),
    .X(_0045_));
 sky130_fd_sc_hd__mux2_1 _2034_ (.A0(_1223_),
    .A1(\simon0.seq[22][1] ),
    .S(_1290_),
    .X(_1292_));
 sky130_fd_sc_hd__clkbuf_1 _2035_ (.A(_1292_),
    .X(_0046_));
 sky130_fd_sc_hd__nor2_1 _2036_ (.A(\simon0.play1.freq[0] ),
    .B(\simon0.play1.tick_counter[0] ),
    .Y(_1293_));
 sky130_fd_sc_hd__and2_1 _2037_ (.A(\simon0.play1.freq[0] ),
    .B(\simon0.play1.tick_counter[0] ),
    .X(_1294_));
 sky130_fd_sc_hd__clkbuf_2 _2038_ (.A(_1294_),
    .X(_1295_));
 sky130_fd_sc_hd__nor3_1 _2039_ (.A(_1201_),
    .B(_1293_),
    .C(_1295_),
    .Y(_0047_));
 sky130_fd_sc_hd__xor2_2 _2040_ (.A(\simon0.play1.freq[1] ),
    .B(\simon0.play1.tick_counter[1] ),
    .X(_1296_));
 sky130_fd_sc_hd__a21oi_1 _2041_ (.A1(_1295_),
    .A2(_1296_),
    .B1(_1123_),
    .Y(_1297_));
 sky130_fd_sc_hd__o21a_1 _2042_ (.A1(_1295_),
    .A2(_1296_),
    .B1(_1297_),
    .X(_0048_));
 sky130_fd_sc_hd__or4_2 _2043_ (.A(\simon0.play1.freq[3] ),
    .B(\simon0.play1.freq[2] ),
    .C(\simon0.play1.freq[1] ),
    .D(\simon0.play1.freq[0] ),
    .X(_1298_));
 sky130_fd_sc_hd__or4_1 _2044_ (.A(\simon0.play1.freq[7] ),
    .B(\simon0.play1.freq[6] ),
    .C(\simon0.play1.freq[5] ),
    .D(\simon0.play1.freq[4] ),
    .X(_1299_));
 sky130_fd_sc_hd__or4_1 _2045_ (.A(\simon0.play1.freq[9] ),
    .B(\simon0.play1.freq[8] ),
    .C(_1298_),
    .D(_1299_),
    .X(_1300_));
 sky130_fd_sc_hd__clkbuf_2 _2046_ (.A(_1300_),
    .X(_1301_));
 sky130_fd_sc_hd__clkbuf_4 _2047_ (.A(_1301_),
    .X(_1302_));
 sky130_fd_sc_hd__clkbuf_4 _2048_ (.A(_1302_),
    .X(_1303_));
 sky130_fd_sc_hd__clkinv_2 _2049_ (.A(net13),
    .Y(_1304_));
 sky130_fd_sc_hd__buf_2 _2050_ (.A(net5),
    .X(_1305_));
 sky130_fd_sc_hd__clkbuf_4 _2051_ (.A(_1305_),
    .X(_1306_));
 sky130_fd_sc_hd__buf_4 _2052_ (.A(_1306_),
    .X(_1307_));
 sky130_fd_sc_hd__nand2_4 _2053_ (.A(_1307_),
    .B(net14),
    .Y(_1308_));
 sky130_fd_sc_hd__nor2_1 _2054_ (.A(_1304_),
    .B(_1308_),
    .Y(_1309_));
 sky130_fd_sc_hd__and3_1 _2055_ (.A(_1306_),
    .B(net10),
    .C(net11),
    .X(_1310_));
 sky130_fd_sc_hd__nand2_1 _2056_ (.A(_1306_),
    .B(net12),
    .Y(_1311_));
 sky130_fd_sc_hd__clkbuf_4 _2057_ (.A(_1311_),
    .X(_1312_));
 sky130_fd_sc_hd__clkbuf_4 _2058_ (.A(net5),
    .X(_1313_));
 sky130_fd_sc_hd__or2b_1 _2059_ (.A(net10),
    .B_N(_1313_),
    .X(_1314_));
 sky130_fd_sc_hd__clkbuf_4 _2060_ (.A(_1314_),
    .X(_1315_));
 sky130_fd_sc_hd__o21bai_2 _2061_ (.A1(net11),
    .A2(_1315_),
    .B1_N(_1310_),
    .Y(_1316_));
 sky130_fd_sc_hd__nor2_1 _2062_ (.A(_1312_),
    .B(_1316_),
    .Y(_1317_));
 sky130_fd_sc_hd__and3_1 _2063_ (.A(_1307_),
    .B(_1304_),
    .C(_1311_),
    .X(_1318_));
 sky130_fd_sc_hd__o21ba_2 _2064_ (.A1(_1304_),
    .A2(_1312_),
    .B1_N(_1318_),
    .X(_1319_));
 sky130_fd_sc_hd__nand2_4 _2065_ (.A(_1306_),
    .B(net11),
    .Y(_1320_));
 sky130_fd_sc_hd__xnor2_1 _2066_ (.A(_1319_),
    .B(_1320_),
    .Y(_1321_));
 sky130_fd_sc_hd__o21a_1 _2067_ (.A1(_1310_),
    .A2(_1317_),
    .B1(_1321_),
    .X(_1322_));
 sky130_fd_sc_hd__nor3_1 _2068_ (.A(_1310_),
    .B(_1317_),
    .C(_1321_),
    .Y(_1323_));
 sky130_fd_sc_hd__or2_1 _2069_ (.A(_1322_),
    .B(_1323_),
    .X(_1324_));
 sky130_fd_sc_hd__nor2_1 _2070_ (.A(_1308_),
    .B(_1324_),
    .Y(_1325_));
 sky130_fd_sc_hd__and2_1 _2071_ (.A(_1308_),
    .B(_1324_),
    .X(_1326_));
 sky130_fd_sc_hd__nor2_1 _2072_ (.A(_1325_),
    .B(_1326_),
    .Y(_1327_));
 sky130_fd_sc_hd__or2b_1 _2073_ (.A(net9),
    .B_N(net5),
    .X(_1328_));
 sky130_fd_sc_hd__clkbuf_4 _2074_ (.A(_1328_),
    .X(_1329_));
 sky130_fd_sc_hd__and2_1 _2075_ (.A(_1315_),
    .B(_1329_),
    .X(_1330_));
 sky130_fd_sc_hd__o21ba_1 _2076_ (.A1(net9),
    .A2(_1315_),
    .B1_N(_1330_),
    .X(_1331_));
 sky130_fd_sc_hd__and3_1 _2077_ (.A(_1307_),
    .B(net11),
    .C(_1331_),
    .X(_1332_));
 sky130_fd_sc_hd__and2_1 _2078_ (.A(_1312_),
    .B(_1316_),
    .X(_1333_));
 sky130_fd_sc_hd__nor2_1 _2079_ (.A(_1317_),
    .B(_1333_),
    .Y(_1334_));
 sky130_fd_sc_hd__o21a_1 _2080_ (.A1(_1330_),
    .A2(_1332_),
    .B1(_1334_),
    .X(_1335_));
 sky130_fd_sc_hd__and2_1 _2081_ (.A(_1307_),
    .B(_1304_),
    .X(_1336_));
 sky130_fd_sc_hd__buf_2 _2082_ (.A(_1336_),
    .X(_1337_));
 sky130_fd_sc_hd__nand2_1 _2083_ (.A(_1337_),
    .B(_1308_),
    .Y(_1338_));
 sky130_fd_sc_hd__o21ai_1 _2084_ (.A1(_1304_),
    .A2(_1308_),
    .B1(_1338_),
    .Y(_1339_));
 sky130_fd_sc_hd__nor3_1 _2085_ (.A(_1334_),
    .B(_1330_),
    .C(_1332_),
    .Y(_1340_));
 sky130_fd_sc_hd__nor2_1 _2086_ (.A(_1335_),
    .B(_1340_),
    .Y(_1341_));
 sky130_fd_sc_hd__and2b_1 _2087_ (.A_N(_1339_),
    .B(_1341_),
    .X(_1342_));
 sky130_fd_sc_hd__nor2_1 _2088_ (.A(_1335_),
    .B(_1342_),
    .Y(_1343_));
 sky130_fd_sc_hd__xnor2_1 _2089_ (.A(_1327_),
    .B(_1343_),
    .Y(_1344_));
 sky130_fd_sc_hd__xnor2_1 _2090_ (.A(_1309_),
    .B(_1344_),
    .Y(_1345_));
 sky130_fd_sc_hd__xor2_1 _2091_ (.A(_1339_),
    .B(_1341_),
    .X(_1346_));
 sky130_fd_sc_hd__xnor2_1 _2092_ (.A(_1320_),
    .B(_1331_),
    .Y(_1347_));
 sky130_fd_sc_hd__a21bo_1 _2093_ (.A1(net23),
    .A2(net9),
    .B1_N(_1305_),
    .X(_1348_));
 sky130_fd_sc_hd__o21ba_1 _2094_ (.A1(net23),
    .A2(_1329_),
    .B1_N(_1348_),
    .X(_1349_));
 sky130_fd_sc_hd__a21oi_1 _2095_ (.A1(_1315_),
    .A2(_1349_),
    .B1(_1348_),
    .Y(_1350_));
 sky130_fd_sc_hd__xnor2_1 _2096_ (.A(_1347_),
    .B(_1350_),
    .Y(_1351_));
 sky130_fd_sc_hd__and2b_1 _2097_ (.A_N(_1350_),
    .B(_1347_),
    .X(_1352_));
 sky130_fd_sc_hd__a21oi_1 _2098_ (.A1(_1319_),
    .A2(_1351_),
    .B1(_1352_),
    .Y(_1353_));
 sky130_fd_sc_hd__xnor2_1 _2099_ (.A(_1346_),
    .B(_1353_),
    .Y(_1354_));
 sky130_fd_sc_hd__or3_1 _2100_ (.A(_1304_),
    .B(_1312_),
    .C(_1354_),
    .X(_1355_));
 sky130_fd_sc_hd__o21ai_1 _2101_ (.A1(_1346_),
    .A2(_1353_),
    .B1(_1355_),
    .Y(_1356_));
 sky130_fd_sc_hd__or2b_1 _2102_ (.A(_1345_),
    .B_N(_1356_),
    .X(_1357_));
 sky130_fd_sc_hd__o21ai_1 _2103_ (.A1(_1304_),
    .A2(_1312_),
    .B1(_1354_),
    .Y(_1358_));
 sky130_fd_sc_hd__nand2_1 _2104_ (.A(_1355_),
    .B(_1358_),
    .Y(_1359_));
 sky130_fd_sc_hd__xnor2_1 _2105_ (.A(_1319_),
    .B(_1351_),
    .Y(_1360_));
 sky130_fd_sc_hd__nor2_1 _2106_ (.A(_1311_),
    .B(_1320_),
    .Y(_1361_));
 sky130_fd_sc_hd__and2_1 _2107_ (.A(_1311_),
    .B(_1320_),
    .X(_1362_));
 sky130_fd_sc_hd__nor2_1 _2108_ (.A(_1361_),
    .B(_1362_),
    .Y(_1363_));
 sky130_fd_sc_hd__xnor2_1 _2109_ (.A(_1315_),
    .B(_1349_),
    .Y(_1364_));
 sky130_fd_sc_hd__inv_2 _2110_ (.A(net22),
    .Y(_1365_));
 sky130_fd_sc_hd__buf_2 _2111_ (.A(net5),
    .X(_1366_));
 sky130_fd_sc_hd__nor2b_4 _2112_ (.A(net23),
    .B_N(_1366_),
    .Y(_1367_));
 sky130_fd_sc_hd__and3_1 _2113_ (.A(_1366_),
    .B(net22),
    .C(net23),
    .X(_1368_));
 sky130_fd_sc_hd__clkbuf_2 _2114_ (.A(_1368_),
    .X(_1369_));
 sky130_fd_sc_hd__a21oi_2 _2115_ (.A1(_1365_),
    .A2(_1367_),
    .B1(_1369_),
    .Y(_1370_));
 sky130_fd_sc_hd__a21oi_1 _2116_ (.A1(_1329_),
    .A2(_1370_),
    .B1(_1369_),
    .Y(_1371_));
 sky130_fd_sc_hd__xor2_1 _2117_ (.A(_1364_),
    .B(_1371_),
    .X(_1372_));
 sky130_fd_sc_hd__nor2_1 _2118_ (.A(_1364_),
    .B(_1371_),
    .Y(_1373_));
 sky130_fd_sc_hd__a21oi_2 _2119_ (.A1(_1363_),
    .A2(_1372_),
    .B1(_1373_),
    .Y(_1374_));
 sky130_fd_sc_hd__xor2_1 _2120_ (.A(_1360_),
    .B(_1374_),
    .X(_1375_));
 sky130_fd_sc_hd__nand2_1 _2121_ (.A(_1361_),
    .B(_1375_),
    .Y(_1376_));
 sky130_fd_sc_hd__o21ai_2 _2122_ (.A1(_1360_),
    .A2(_1374_),
    .B1(_1376_),
    .Y(_1377_));
 sky130_fd_sc_hd__or2b_1 _2123_ (.A(_1359_),
    .B_N(_1377_),
    .X(_1378_));
 sky130_fd_sc_hd__xor2_1 _2124_ (.A(_1345_),
    .B(_1356_),
    .X(_1379_));
 sky130_fd_sc_hd__nor2_1 _2125_ (.A(_1378_),
    .B(_1379_),
    .Y(_1380_));
 sky130_fd_sc_hd__and2_1 _2126_ (.A(_1378_),
    .B(_1379_),
    .X(_1381_));
 sky130_fd_sc_hd__nor2_1 _2127_ (.A(_1380_),
    .B(_1381_),
    .Y(_1382_));
 sky130_fd_sc_hd__and3_1 _2128_ (.A(_1305_),
    .B(net21),
    .C(net22),
    .X(_1383_));
 sky130_fd_sc_hd__o21ai_1 _2129_ (.A1(net21),
    .A2(net22),
    .B1(_1313_),
    .Y(_1384_));
 sky130_fd_sc_hd__or3_1 _2130_ (.A(_1367_),
    .B(_1383_),
    .C(_1384_),
    .X(_1385_));
 sky130_fd_sc_hd__nand2b_1 _2131_ (.A_N(_1383_),
    .B(_1385_),
    .Y(_1386_));
 sky130_fd_sc_hd__xor2_1 _2132_ (.A(_1329_),
    .B(_1370_),
    .X(_1387_));
 sky130_fd_sc_hd__nor2_1 _2133_ (.A(_1386_),
    .B(_1387_),
    .Y(_1388_));
 sky130_fd_sc_hd__nand2_1 _2134_ (.A(_1386_),
    .B(_1387_),
    .Y(_1389_));
 sky130_fd_sc_hd__o21a_1 _2135_ (.A1(_1316_),
    .A2(_1388_),
    .B1(_1389_),
    .X(_1390_));
 sky130_fd_sc_hd__xnor2_1 _2136_ (.A(_1363_),
    .B(_1372_),
    .Y(_1391_));
 sky130_fd_sc_hd__xor2_1 _2137_ (.A(_1390_),
    .B(_1391_),
    .X(_1392_));
 sky130_fd_sc_hd__xnor2_1 _2138_ (.A(_1310_),
    .B(_1392_),
    .Y(_1393_));
 sky130_fd_sc_hd__o21ai_1 _2139_ (.A1(_1383_),
    .A2(_1384_),
    .B1(_1367_),
    .Y(_1394_));
 sky130_fd_sc_hd__nand2_2 _2140_ (.A(_1313_),
    .B(net22),
    .Y(_1395_));
 sky130_fd_sc_hd__o21ai_1 _2141_ (.A1(net20),
    .A2(net21),
    .B1(_1313_),
    .Y(_1396_));
 sky130_fd_sc_hd__and3_1 _2142_ (.A(_1305_),
    .B(net20),
    .C(net21),
    .X(_1397_));
 sky130_fd_sc_hd__o21bai_1 _2143_ (.A1(_1395_),
    .A2(_1396_),
    .B1_N(_1397_),
    .Y(_1398_));
 sky130_fd_sc_hd__a21o_1 _2144_ (.A1(_1385_),
    .A2(_1394_),
    .B1(_1398_),
    .X(_1399_));
 sky130_fd_sc_hd__and3_1 _2145_ (.A(_1385_),
    .B(_1398_),
    .C(_1394_),
    .X(_1400_));
 sky130_fd_sc_hd__a21oi_1 _2146_ (.A1(_1331_),
    .A2(_1399_),
    .B1(_1400_),
    .Y(_1401_));
 sky130_fd_sc_hd__xor2_1 _2147_ (.A(_1386_),
    .B(_1387_),
    .X(_1402_));
 sky130_fd_sc_hd__xnor2_1 _2148_ (.A(_1316_),
    .B(_1402_),
    .Y(_1403_));
 sky130_fd_sc_hd__xnor2_1 _2149_ (.A(_1401_),
    .B(_1403_),
    .Y(_1404_));
 sky130_fd_sc_hd__and2b_1 _2150_ (.A_N(_1401_),
    .B(_1403_),
    .X(_1405_));
 sky130_fd_sc_hd__a21o_1 _2151_ (.A1(_1330_),
    .A2(_1404_),
    .B1(_1405_),
    .X(_1406_));
 sky130_fd_sc_hd__or2b_1 _2152_ (.A(_1393_),
    .B_N(_1406_),
    .X(_1407_));
 sky130_fd_sc_hd__and2_1 _2153_ (.A(_1307_),
    .B(net14),
    .X(_1408_));
 sky130_fd_sc_hd__xnor2_1 _2154_ (.A(_1406_),
    .B(_1393_),
    .Y(_1409_));
 sky130_fd_sc_hd__nand2_1 _2155_ (.A(_1408_),
    .B(_1409_),
    .Y(_1410_));
 sky130_fd_sc_hd__or2_1 _2156_ (.A(_1361_),
    .B(_1375_),
    .X(_1411_));
 sky130_fd_sc_hd__nand2_1 _2157_ (.A(_1376_),
    .B(_1411_),
    .Y(_1412_));
 sky130_fd_sc_hd__nor2_1 _2158_ (.A(_1390_),
    .B(_1391_),
    .Y(_1413_));
 sky130_fd_sc_hd__a21o_1 _2159_ (.A1(_1310_),
    .A2(_1392_),
    .B1(_1413_),
    .X(_1414_));
 sky130_fd_sc_hd__xor2_1 _2160_ (.A(_1412_),
    .B(_1414_),
    .X(_1415_));
 sky130_fd_sc_hd__a21oi_2 _2161_ (.A1(_1407_),
    .A2(_1410_),
    .B1(_1415_),
    .Y(_1416_));
 sky130_fd_sc_hd__and3_1 _2162_ (.A(_1415_),
    .B(_1407_),
    .C(_1410_),
    .X(_1417_));
 sky130_fd_sc_hd__nor2_2 _2163_ (.A(_1416_),
    .B(_1417_),
    .Y(_1418_));
 sky130_fd_sc_hd__nor2_1 _2164_ (.A(_1383_),
    .B(_1384_),
    .Y(_1419_));
 sky130_fd_sc_hd__nand2_2 _2165_ (.A(_1313_),
    .B(net20),
    .Y(_1420_));
 sky130_fd_sc_hd__and3_1 _2166_ (.A(_1313_),
    .B(net18),
    .C(net19),
    .X(_1421_));
 sky130_fd_sc_hd__or3b_1 _2167_ (.A(net18),
    .B(net19),
    .C_N(_1305_),
    .X(_1422_));
 sky130_fd_sc_hd__or3b_1 _2168_ (.A(_1420_),
    .B(_1421_),
    .C_N(_1422_),
    .X(_1423_));
 sky130_fd_sc_hd__nand3_2 _2169_ (.A(_1313_),
    .B(net18),
    .C(net19),
    .Y(_1424_));
 sky130_fd_sc_hd__a21bo_1 _2170_ (.A1(_1424_),
    .A2(_1422_),
    .B1_N(_1420_),
    .X(_1425_));
 sky130_fd_sc_hd__or2b_1 _2171_ (.A(net19),
    .B_N(_1305_),
    .X(_1426_));
 sky130_fd_sc_hd__o21a_1 _2172_ (.A1(net17),
    .A2(net18),
    .B1(_1366_),
    .X(_1427_));
 sky130_fd_sc_hd__and3_1 _2173_ (.A(_1366_),
    .B(net17),
    .C(net18),
    .X(_1428_));
 sky130_fd_sc_hd__a21o_1 _2174_ (.A1(_1426_),
    .A2(_1427_),
    .B1(_1428_),
    .X(_1429_));
 sky130_fd_sc_hd__a21o_1 _2175_ (.A1(_1423_),
    .A2(_1425_),
    .B1(_1429_),
    .X(_1430_));
 sky130_fd_sc_hd__nand3_1 _2176_ (.A(_1429_),
    .B(_1423_),
    .C(_1425_),
    .Y(_1431_));
 sky130_fd_sc_hd__a21bo_1 _2177_ (.A1(_1419_),
    .A2(_1430_),
    .B1_N(_1431_),
    .X(_1432_));
 sky130_fd_sc_hd__a31o_1 _2178_ (.A1(_1307_),
    .A2(net20),
    .A3(_1422_),
    .B1(_1421_),
    .X(_1433_));
 sky130_fd_sc_hd__nand2_2 _2179_ (.A(_1306_),
    .B(net21),
    .Y(_1434_));
 sky130_fd_sc_hd__and3_1 _2180_ (.A(_1313_),
    .B(net19),
    .C(net20),
    .X(_1435_));
 sky130_fd_sc_hd__or3b_1 _2181_ (.A(net19),
    .B(net20),
    .C_N(_1305_),
    .X(_1436_));
 sky130_fd_sc_hd__or3b_1 _2182_ (.A(_1434_),
    .B(_1435_),
    .C_N(_1436_),
    .X(_1437_));
 sky130_fd_sc_hd__nand3_1 _2183_ (.A(_1306_),
    .B(net19),
    .C(net20),
    .Y(_1438_));
 sky130_fd_sc_hd__a21bo_1 _2184_ (.A1(_1438_),
    .A2(_1436_),
    .B1_N(_1434_),
    .X(_1439_));
 sky130_fd_sc_hd__nand3_1 _2185_ (.A(_1433_),
    .B(_1437_),
    .C(_1439_),
    .Y(_1440_));
 sky130_fd_sc_hd__a21o_1 _2186_ (.A1(_1437_),
    .A2(_1439_),
    .B1(_1433_),
    .X(_1441_));
 sky130_fd_sc_hd__nand3_1 _2187_ (.A(_1370_),
    .B(_1440_),
    .C(_1441_),
    .Y(_1442_));
 sky130_fd_sc_hd__a21o_1 _2188_ (.A1(_1440_),
    .A2(_1441_),
    .B1(_1370_),
    .X(_1443_));
 sky130_fd_sc_hd__nand3_1 _2189_ (.A(_1432_),
    .B(_1442_),
    .C(_1443_),
    .Y(_1444_));
 sky130_fd_sc_hd__a21o_1 _2190_ (.A1(_1442_),
    .A2(_1443_),
    .B1(_1432_),
    .X(_1445_));
 sky130_fd_sc_hd__nand3_1 _2191_ (.A(_1383_),
    .B(_1444_),
    .C(_1445_),
    .Y(_1446_));
 sky130_fd_sc_hd__nand3_1 _2192_ (.A(_1419_),
    .B(_1431_),
    .C(_1430_),
    .Y(_1447_));
 sky130_fd_sc_hd__a21o_1 _2193_ (.A1(_1431_),
    .A2(_1430_),
    .B1(_1419_),
    .X(_1448_));
 sky130_fd_sc_hd__nor2_1 _2194_ (.A(_1397_),
    .B(_1396_),
    .Y(_1449_));
 sky130_fd_sc_hd__and2b_1 _2195_ (.A_N(net19),
    .B(_1366_),
    .X(_1450_));
 sky130_fd_sc_hd__or3b_1 _2196_ (.A(_1428_),
    .B(_1450_),
    .C_N(_1427_),
    .X(_1451_));
 sky130_fd_sc_hd__nand3_2 _2197_ (.A(_1305_),
    .B(net17),
    .C(net18),
    .Y(_1452_));
 sky130_fd_sc_hd__a21o_1 _2198_ (.A1(_1452_),
    .A2(_1427_),
    .B1(_1426_),
    .X(_1453_));
 sky130_fd_sc_hd__o21a_1 _2199_ (.A1(net16),
    .A2(net17),
    .B1(_1366_),
    .X(_0172_));
 sky130_fd_sc_hd__and3_1 _2200_ (.A(_1366_),
    .B(net16),
    .C(net17),
    .X(_0173_));
 sky130_fd_sc_hd__a31o_1 _2201_ (.A1(_1313_),
    .A2(net18),
    .A3(_0172_),
    .B1(_0173_),
    .X(_0174_));
 sky130_fd_sc_hd__a21o_1 _2202_ (.A1(_1451_),
    .A2(_1453_),
    .B1(_0174_),
    .X(_0175_));
 sky130_fd_sc_hd__nand3_1 _2203_ (.A(_1451_),
    .B(_0174_),
    .C(_1453_),
    .Y(_0176_));
 sky130_fd_sc_hd__a21bo_1 _2204_ (.A1(_1449_),
    .A2(_0175_),
    .B1_N(_0176_),
    .X(_0177_));
 sky130_fd_sc_hd__a21o_1 _2205_ (.A1(_1447_),
    .A2(_1448_),
    .B1(_0177_),
    .X(_0178_));
 sky130_fd_sc_hd__nand3_1 _2206_ (.A(_1447_),
    .B(_0177_),
    .C(_1448_),
    .Y(_0179_));
 sky130_fd_sc_hd__a21bo_1 _2207_ (.A1(_1397_),
    .A2(_0178_),
    .B1_N(_0179_),
    .X(_0180_));
 sky130_fd_sc_hd__a21o_1 _2208_ (.A1(_1444_),
    .A2(_1445_),
    .B1(_1383_),
    .X(_0181_));
 sky130_fd_sc_hd__nand3_1 _2209_ (.A(_1446_),
    .B(_0180_),
    .C(_0181_),
    .Y(_0182_));
 sky130_fd_sc_hd__a21o_1 _2210_ (.A1(_1446_),
    .A2(_0181_),
    .B1(_0180_),
    .X(_0183_));
 sky130_fd_sc_hd__nand3_1 _2211_ (.A(_1315_),
    .B(_0182_),
    .C(_0183_),
    .Y(_0184_));
 sky130_fd_sc_hd__a21o_1 _2212_ (.A1(_0182_),
    .A2(_0183_),
    .B1(_1315_),
    .X(_0185_));
 sky130_fd_sc_hd__nand3_1 _2213_ (.A(_1397_),
    .B(_0179_),
    .C(_0178_),
    .Y(_0186_));
 sky130_fd_sc_hd__a21o_1 _2214_ (.A1(_0179_),
    .A2(_0178_),
    .B1(_1397_),
    .X(_0187_));
 sky130_fd_sc_hd__nand3_1 _2215_ (.A(_1449_),
    .B(_0176_),
    .C(_0175_),
    .Y(_0188_));
 sky130_fd_sc_hd__a21o_1 _2216_ (.A1(_0176_),
    .A2(_0175_),
    .B1(_1449_),
    .X(_0189_));
 sky130_fd_sc_hd__and2_1 _2217_ (.A(_1438_),
    .B(_1436_),
    .X(_0190_));
 sky130_fd_sc_hd__nand2_2 _2218_ (.A(_1366_),
    .B(net18),
    .Y(_0191_));
 sky130_fd_sc_hd__or3b_1 _2219_ (.A(_0191_),
    .B(_0173_),
    .C_N(_0172_),
    .X(_0192_));
 sky130_fd_sc_hd__nand3_2 _2220_ (.A(_1305_),
    .B(net16),
    .C(net17),
    .Y(_0193_));
 sky130_fd_sc_hd__a21bo_1 _2221_ (.A1(_0193_),
    .A2(_0172_),
    .B1_N(_0191_),
    .X(_0194_));
 sky130_fd_sc_hd__nand2_2 _2222_ (.A(net5),
    .B(net17),
    .Y(_0195_));
 sky130_fd_sc_hd__o21ai_1 _2223_ (.A1(net15),
    .A2(net16),
    .B1(_1366_),
    .Y(_0196_));
 sky130_fd_sc_hd__and3_1 _2224_ (.A(net5),
    .B(net15),
    .C(net16),
    .X(_0197_));
 sky130_fd_sc_hd__o21bai_1 _2225_ (.A1(_0195_),
    .A2(_0196_),
    .B1_N(_0197_),
    .Y(_0198_));
 sky130_fd_sc_hd__a21o_1 _2226_ (.A1(_0192_),
    .A2(_0194_),
    .B1(_0198_),
    .X(_0199_));
 sky130_fd_sc_hd__nand3_1 _2227_ (.A(_0192_),
    .B(_0198_),
    .C(_0194_),
    .Y(_0200_));
 sky130_fd_sc_hd__a21bo_1 _2228_ (.A1(_0190_),
    .A2(_0199_),
    .B1_N(_0200_),
    .X(_0201_));
 sky130_fd_sc_hd__a21oi_1 _2229_ (.A1(_0188_),
    .A2(_0189_),
    .B1(_0201_),
    .Y(_0202_));
 sky130_fd_sc_hd__and3_1 _2230_ (.A(_0188_),
    .B(_0201_),
    .C(_0189_),
    .X(_0203_));
 sky130_fd_sc_hd__o21bai_1 _2231_ (.A1(_1438_),
    .A2(_0202_),
    .B1_N(_0203_),
    .Y(_0204_));
 sky130_fd_sc_hd__a21o_1 _2232_ (.A1(_0186_),
    .A2(_0187_),
    .B1(_0204_),
    .X(_0205_));
 sky130_fd_sc_hd__and3_1 _2233_ (.A(_0186_),
    .B(_0204_),
    .C(_0187_),
    .X(_0206_));
 sky130_fd_sc_hd__a21o_1 _2234_ (.A1(_1329_),
    .A2(_0205_),
    .B1(_0206_),
    .X(_0207_));
 sky130_fd_sc_hd__a21oi_1 _2235_ (.A1(_0184_),
    .A2(_0185_),
    .B1(_0207_),
    .Y(_0208_));
 sky130_fd_sc_hd__and2b_1 _2236_ (.A_N(_0206_),
    .B(_0205_),
    .X(_0209_));
 sky130_fd_sc_hd__xor2_2 _2237_ (.A(_1329_),
    .B(_0209_),
    .X(_0210_));
 sky130_fd_sc_hd__or3_1 _2238_ (.A(_1438_),
    .B(_0203_),
    .C(_0202_),
    .X(_0211_));
 sky130_fd_sc_hd__nand3_1 _2239_ (.A(_0190_),
    .B(_0200_),
    .C(_0199_),
    .Y(_0212_));
 sky130_fd_sc_hd__a21o_1 _2240_ (.A1(_0200_),
    .A2(_0199_),
    .B1(_0190_),
    .X(_0213_));
 sky130_fd_sc_hd__and2_1 _2241_ (.A(_1424_),
    .B(_1422_),
    .X(_0214_));
 sky130_fd_sc_hd__or3_1 _2242_ (.A(_0195_),
    .B(_0197_),
    .C(_0196_),
    .X(_0215_));
 sky130_fd_sc_hd__o21ai_1 _2243_ (.A1(_0197_),
    .A2(_0196_),
    .B1(_0195_),
    .Y(_0216_));
 sky130_fd_sc_hd__and3_1 _2244_ (.A(net5),
    .B(net8),
    .C(net15),
    .X(_0217_));
 sky130_fd_sc_hd__o211a_1 _2245_ (.A1(net8),
    .A2(net15),
    .B1(net16),
    .C1(_1366_),
    .X(_0218_));
 sky130_fd_sc_hd__or2_1 _2246_ (.A(_0217_),
    .B(_0218_),
    .X(_0219_));
 sky130_fd_sc_hd__a21o_1 _2247_ (.A1(_0215_),
    .A2(_0216_),
    .B1(_0219_),
    .X(_0220_));
 sky130_fd_sc_hd__nand3_1 _2248_ (.A(_0215_),
    .B(_0216_),
    .C(_0219_),
    .Y(_0221_));
 sky130_fd_sc_hd__a21bo_1 _2249_ (.A1(_0214_),
    .A2(_0220_),
    .B1_N(_0221_),
    .X(_0222_));
 sky130_fd_sc_hd__a21oi_1 _2250_ (.A1(_0212_),
    .A2(_0213_),
    .B1(_0222_),
    .Y(_0223_));
 sky130_fd_sc_hd__and3_1 _2251_ (.A(_0212_),
    .B(_0222_),
    .C(_0213_),
    .X(_0224_));
 sky130_fd_sc_hd__o21bai_1 _2252_ (.A1(_1424_),
    .A2(_0223_),
    .B1_N(_0224_),
    .Y(_0225_));
 sky130_fd_sc_hd__o21ai_1 _2253_ (.A1(_0203_),
    .A2(_0202_),
    .B1(_1438_),
    .Y(_0226_));
 sky130_fd_sc_hd__and3_1 _2254_ (.A(_0211_),
    .B(_0225_),
    .C(_0226_),
    .X(_0227_));
 sky130_fd_sc_hd__a21oi_1 _2255_ (.A1(_0211_),
    .A2(_0226_),
    .B1(_0225_),
    .Y(_0228_));
 sky130_fd_sc_hd__or3_1 _2256_ (.A(_1367_),
    .B(_0227_),
    .C(_0228_),
    .X(_0229_));
 sky130_fd_sc_hd__or2b_1 _2257_ (.A(_0227_),
    .B_N(_0229_),
    .X(_0230_));
 sky130_fd_sc_hd__nand2_1 _2258_ (.A(_0210_),
    .B(_0230_),
    .Y(_0231_));
 sky130_fd_sc_hd__and3_1 _2259_ (.A(_0184_),
    .B(_0185_),
    .C(_0207_),
    .X(_0232_));
 sky130_fd_sc_hd__o21ba_1 _2260_ (.A1(_0208_),
    .A2(_0231_),
    .B1_N(_0232_),
    .X(_0233_));
 sky130_fd_sc_hd__xor2_2 _2261_ (.A(_0210_),
    .B(_0230_),
    .X(_0234_));
 sky130_fd_sc_hd__and2_1 _2262_ (.A(_1307_),
    .B(net22),
    .X(_0235_));
 sky130_fd_sc_hd__or3_1 _2263_ (.A(_1424_),
    .B(_0224_),
    .C(_0223_),
    .X(_0236_));
 sky130_fd_sc_hd__nand3_1 _2264_ (.A(_0214_),
    .B(_0221_),
    .C(_0220_),
    .Y(_0237_));
 sky130_fd_sc_hd__a21o_1 _2265_ (.A1(_0221_),
    .A2(_0220_),
    .B1(_0214_),
    .X(_0238_));
 sky130_fd_sc_hd__nand2_1 _2266_ (.A(_1452_),
    .B(_1427_),
    .Y(_0239_));
 sky130_fd_sc_hd__o31ai_1 _2267_ (.A1(net8),
    .A2(net15),
    .A3(net16),
    .B1(_1305_),
    .Y(_0240_));
 sky130_fd_sc_hd__or2_2 _2268_ (.A(_0218_),
    .B(_0240_),
    .X(_0241_));
 sky130_fd_sc_hd__nand2_2 _2269_ (.A(_1313_),
    .B(net8),
    .Y(_0242_));
 sky130_fd_sc_hd__nand2_1 _2270_ (.A(_1306_),
    .B(net16),
    .Y(_0243_));
 sky130_fd_sc_hd__nor2_1 _2271_ (.A(_0242_),
    .B(_0243_),
    .Y(_0244_));
 sky130_fd_sc_hd__and2_1 _2272_ (.A(_1306_),
    .B(net15),
    .X(_0245_));
 sky130_fd_sc_hd__a2bb2o_1 _2273_ (.A1_N(_0239_),
    .A2_N(_0241_),
    .B1(_0244_),
    .B2(_0245_),
    .X(_0246_));
 sky130_fd_sc_hd__a21oi_1 _2274_ (.A1(_0237_),
    .A2(_0238_),
    .B1(_0246_),
    .Y(_0247_));
 sky130_fd_sc_hd__and3_1 _2275_ (.A(_0237_),
    .B(_0238_),
    .C(_0246_),
    .X(_0248_));
 sky130_fd_sc_hd__o21bai_1 _2276_ (.A1(_1452_),
    .A2(_0247_),
    .B1_N(_0248_),
    .Y(_0249_));
 sky130_fd_sc_hd__o21ai_1 _2277_ (.A1(_0224_),
    .A2(_0223_),
    .B1(_1424_),
    .Y(_0250_));
 sky130_fd_sc_hd__nand3_1 _2278_ (.A(_0236_),
    .B(_0249_),
    .C(_0250_),
    .Y(_0251_));
 sky130_fd_sc_hd__a21o_1 _2279_ (.A1(_0236_),
    .A2(_0250_),
    .B1(_0249_),
    .X(_0252_));
 sky130_fd_sc_hd__nand3_1 _2280_ (.A(_0235_),
    .B(_0251_),
    .C(_0252_),
    .Y(_0253_));
 sky130_fd_sc_hd__a21o_1 _2281_ (.A1(_0251_),
    .A2(_0252_),
    .B1(_0235_),
    .X(_0254_));
 sky130_fd_sc_hd__or3_1 _2282_ (.A(_1452_),
    .B(_0248_),
    .C(_0247_),
    .X(_0255_));
 sky130_fd_sc_hd__o21ai_1 _2283_ (.A1(_0248_),
    .A2(_0247_),
    .B1(_1452_),
    .Y(_0256_));
 sky130_fd_sc_hd__xnor2_1 _2284_ (.A(_0239_),
    .B(_0241_),
    .Y(_0257_));
 sky130_fd_sc_hd__nand2_1 _2285_ (.A(_0193_),
    .B(_0172_),
    .Y(_0258_));
 sky130_fd_sc_hd__o21ai_1 _2286_ (.A1(net8),
    .A2(net15),
    .B1(_1306_),
    .Y(_0259_));
 sky130_fd_sc_hd__or3_1 _2287_ (.A(_0258_),
    .B(_0217_),
    .C(_0259_),
    .X(_0260_));
 sky130_fd_sc_hd__xor2_1 _2288_ (.A(_0191_),
    .B(_0241_),
    .X(_0261_));
 sky130_fd_sc_hd__nor2_1 _2289_ (.A(_0193_),
    .B(_0261_),
    .Y(_0262_));
 sky130_fd_sc_hd__o21bai_1 _2290_ (.A1(_0257_),
    .A2(_0260_),
    .B1_N(_0262_),
    .Y(_0263_));
 sky130_fd_sc_hd__a21oi_1 _2291_ (.A1(_0255_),
    .A2(_0256_),
    .B1(_0263_),
    .Y(_0264_));
 sky130_fd_sc_hd__and3_1 _2292_ (.A(_0255_),
    .B(_0263_),
    .C(_0256_),
    .X(_0265_));
 sky130_fd_sc_hd__o21bai_1 _2293_ (.A1(_1434_),
    .A2(_0264_),
    .B1_N(_0265_),
    .Y(_0266_));
 sky130_fd_sc_hd__nand3_1 _2294_ (.A(_0253_),
    .B(_0254_),
    .C(_0266_),
    .Y(_0267_));
 sky130_fd_sc_hd__o21ai_1 _2295_ (.A1(_0227_),
    .A2(_0228_),
    .B1(_1367_),
    .Y(_0268_));
 sky130_fd_sc_hd__a21bo_1 _2296_ (.A1(_0235_),
    .A2(_0252_),
    .B1_N(_0251_),
    .X(_0269_));
 sky130_fd_sc_hd__nand3_1 _2297_ (.A(_0229_),
    .B(_0268_),
    .C(_0269_),
    .Y(_0270_));
 sky130_fd_sc_hd__a21oi_1 _2298_ (.A1(_0229_),
    .A2(_0268_),
    .B1(_0269_),
    .Y(_0271_));
 sky130_fd_sc_hd__a21oi_1 _2299_ (.A1(_0267_),
    .A2(_0270_),
    .B1(_0271_),
    .Y(_0272_));
 sky130_fd_sc_hd__nor2_1 _2300_ (.A(_0232_),
    .B(_0208_),
    .Y(_0273_));
 sky130_fd_sc_hd__nand3_1 _2301_ (.A(_0234_),
    .B(_0272_),
    .C(_0273_),
    .Y(_0274_));
 sky130_fd_sc_hd__nor3_1 _2302_ (.A(_1434_),
    .B(_0265_),
    .C(_0264_),
    .Y(_0275_));
 sky130_fd_sc_hd__o21a_1 _2303_ (.A1(_0265_),
    .A2(_0264_),
    .B1(_1434_),
    .X(_0276_));
 sky130_fd_sc_hd__xnor2_1 _2304_ (.A(_0257_),
    .B(_0260_),
    .Y(_0277_));
 sky130_fd_sc_hd__a21o_1 _2305_ (.A1(_0193_),
    .A2(_0277_),
    .B1(_0262_),
    .X(_0278_));
 sky130_fd_sc_hd__o21ai_1 _2306_ (.A1(_0217_),
    .A2(_0259_),
    .B1(_0258_),
    .Y(_0279_));
 sky130_fd_sc_hd__nand3_1 _2307_ (.A(_0219_),
    .B(_0260_),
    .C(_0279_),
    .Y(_0280_));
 sky130_fd_sc_hd__xnor2_1 _2308_ (.A(_0278_),
    .B(_0280_),
    .Y(_0281_));
 sky130_fd_sc_hd__or2_1 _2309_ (.A(_0278_),
    .B(_0280_),
    .X(_0282_));
 sky130_fd_sc_hd__o21ai_1 _2310_ (.A1(_1420_),
    .A2(_0281_),
    .B1(_0282_),
    .Y(_0283_));
 sky130_fd_sc_hd__inv_2 _2311_ (.A(_0283_),
    .Y(_0284_));
 sky130_fd_sc_hd__o21ai_1 _2312_ (.A1(_0275_),
    .A2(_0276_),
    .B1(_0284_),
    .Y(_0285_));
 sky130_fd_sc_hd__xnor2_2 _2313_ (.A(_1420_),
    .B(_0281_),
    .Y(_0286_));
 sky130_fd_sc_hd__xnor2_1 _2314_ (.A(_0195_),
    .B(_0240_),
    .Y(_0287_));
 sky130_fd_sc_hd__o2bb2a_1 _2315_ (.A1_N(_0173_),
    .A2_N(_0217_),
    .B1(_0287_),
    .B2(_1450_),
    .X(_0288_));
 sky130_fd_sc_hd__xor2_2 _2316_ (.A(_0286_),
    .B(_0288_),
    .X(_0289_));
 sky130_fd_sc_hd__xnor2_2 _2317_ (.A(_1450_),
    .B(_0287_),
    .Y(_0290_));
 sky130_fd_sc_hd__nor3_1 _2318_ (.A(_0195_),
    .B(_0217_),
    .C(_0259_),
    .Y(_0291_));
 sky130_fd_sc_hd__o21a_1 _2319_ (.A1(_0217_),
    .A2(_0259_),
    .B1(_0195_),
    .X(_0292_));
 sky130_fd_sc_hd__nor2_1 _2320_ (.A(_0291_),
    .B(_0292_),
    .Y(_0293_));
 sky130_fd_sc_hd__and2_1 _2321_ (.A(_0244_),
    .B(_0293_),
    .X(_0294_));
 sky130_fd_sc_hd__o21ai_1 _2322_ (.A1(_0291_),
    .A2(_0294_),
    .B1(_0261_),
    .Y(_0295_));
 sky130_fd_sc_hd__o21a_1 _2323_ (.A1(_0191_),
    .A2(_0241_),
    .B1(_0295_),
    .X(_0296_));
 sky130_fd_sc_hd__nor2_1 _2324_ (.A(_0290_),
    .B(_0296_),
    .Y(_0297_));
 sky130_fd_sc_hd__nor2_1 _2325_ (.A(_0286_),
    .B(_0288_),
    .Y(_0298_));
 sky130_fd_sc_hd__a21o_1 _2326_ (.A1(_0289_),
    .A2(_0297_),
    .B1(_0298_),
    .X(_0299_));
 sky130_fd_sc_hd__or3_1 _2327_ (.A(_0275_),
    .B(_0276_),
    .C(_0284_),
    .X(_0300_));
 sky130_fd_sc_hd__a21bo_1 _2328_ (.A1(_0285_),
    .A2(_0299_),
    .B1_N(_0300_),
    .X(_0301_));
 sky130_fd_sc_hd__a21o_1 _2329_ (.A1(_0253_),
    .A2(_0254_),
    .B1(_0266_),
    .X(_0302_));
 sky130_fd_sc_hd__and4b_1 _2330_ (.A_N(_0271_),
    .B(_0267_),
    .C(_0270_),
    .D(_0302_),
    .X(_0303_));
 sky130_fd_sc_hd__nand4_1 _2331_ (.A(_0234_),
    .B(_0301_),
    .C(_0303_),
    .D(_0273_),
    .Y(_0304_));
 sky130_fd_sc_hd__nand2_1 _2332_ (.A(_1444_),
    .B(_1446_),
    .Y(_0305_));
 sky130_fd_sc_hd__and2_1 _2333_ (.A(_1440_),
    .B(_1442_),
    .X(_0306_));
 sky130_fd_sc_hd__or3_1 _2334_ (.A(_1395_),
    .B(_1397_),
    .C(_1396_),
    .X(_0307_));
 sky130_fd_sc_hd__a31o_1 _2335_ (.A1(_1306_),
    .A2(net21),
    .A3(_1436_),
    .B1(_1435_),
    .X(_0308_));
 sky130_fd_sc_hd__o21ai_1 _2336_ (.A1(_1397_),
    .A2(_1396_),
    .B1(_1395_),
    .Y(_0309_));
 sky130_fd_sc_hd__and3_1 _2337_ (.A(_0307_),
    .B(_0308_),
    .C(_0309_),
    .X(_0310_));
 sky130_fd_sc_hd__a21o_1 _2338_ (.A1(_0307_),
    .A2(_0309_),
    .B1(_0308_),
    .X(_0311_));
 sky130_fd_sc_hd__and2b_1 _2339_ (.A_N(_0310_),
    .B(_0311_),
    .X(_0312_));
 sky130_fd_sc_hd__xnor2_1 _2340_ (.A(_1349_),
    .B(_0312_),
    .Y(_0313_));
 sky130_fd_sc_hd__xor2_1 _2341_ (.A(_0306_),
    .B(_0313_),
    .X(_0314_));
 sky130_fd_sc_hd__xnor2_1 _2342_ (.A(_1369_),
    .B(_0314_),
    .Y(_0315_));
 sky130_fd_sc_hd__xor2_1 _2343_ (.A(_0305_),
    .B(_0315_),
    .X(_0316_));
 sky130_fd_sc_hd__xnor2_1 _2344_ (.A(_1320_),
    .B(_0316_),
    .Y(_0317_));
 sky130_fd_sc_hd__nand2_1 _2345_ (.A(_0182_),
    .B(_0184_),
    .Y(_0318_));
 sky130_fd_sc_hd__xor2_1 _2346_ (.A(_0317_),
    .B(_0318_),
    .X(_0319_));
 sky130_fd_sc_hd__a31o_2 _2347_ (.A1(_0233_),
    .A2(_0274_),
    .A3(_0304_),
    .B1(_0319_),
    .X(_0320_));
 sky130_fd_sc_hd__or2b_1 _2348_ (.A(_0315_),
    .B_N(_0305_),
    .X(_0321_));
 sky130_fd_sc_hd__or2_1 _2349_ (.A(_1320_),
    .B(_0316_),
    .X(_0322_));
 sky130_fd_sc_hd__nor2_1 _2350_ (.A(_0306_),
    .B(_0313_),
    .Y(_0323_));
 sky130_fd_sc_hd__a21oi_1 _2351_ (.A1(_1369_),
    .A2(_0314_),
    .B1(_0323_),
    .Y(_0324_));
 sky130_fd_sc_hd__a21o_1 _2352_ (.A1(_1349_),
    .A2(_0311_),
    .B1(_0310_),
    .X(_0325_));
 sky130_fd_sc_hd__or2b_1 _2353_ (.A(_1400_),
    .B_N(_1399_),
    .X(_0326_));
 sky130_fd_sc_hd__xnor2_1 _2354_ (.A(_1331_),
    .B(_0326_),
    .Y(_0327_));
 sky130_fd_sc_hd__xor2_1 _2355_ (.A(_0325_),
    .B(_0327_),
    .X(_0328_));
 sky130_fd_sc_hd__xnor2_1 _2356_ (.A(_1348_),
    .B(_0328_),
    .Y(_0329_));
 sky130_fd_sc_hd__xnor2_1 _2357_ (.A(_0324_),
    .B(_0329_),
    .Y(_0330_));
 sky130_fd_sc_hd__xnor2_1 _2358_ (.A(_1312_),
    .B(_0330_),
    .Y(_0331_));
 sky130_fd_sc_hd__and3_1 _2359_ (.A(_0321_),
    .B(_0322_),
    .C(_0331_),
    .X(_0332_));
 sky130_fd_sc_hd__a21o_1 _2360_ (.A1(_0321_),
    .A2(_0322_),
    .B1(_0331_),
    .X(_0333_));
 sky130_fd_sc_hd__or2b_2 _2361_ (.A(_0332_),
    .B_N(_0333_),
    .X(_0334_));
 sky130_fd_sc_hd__xnor2_1 _2362_ (.A(_1308_),
    .B(_1409_),
    .Y(_0335_));
 sky130_fd_sc_hd__and2_1 _2363_ (.A(_0325_),
    .B(_0327_),
    .X(_0336_));
 sky130_fd_sc_hd__a21oi_1 _2364_ (.A1(_1348_),
    .A2(_0328_),
    .B1(_0336_),
    .Y(_0337_));
 sky130_fd_sc_hd__xnor2_1 _2365_ (.A(_1330_),
    .B(_1404_),
    .Y(_0338_));
 sky130_fd_sc_hd__xnor2_1 _2366_ (.A(_0337_),
    .B(_0338_),
    .Y(_0339_));
 sky130_fd_sc_hd__or2_1 _2367_ (.A(_0337_),
    .B(_0338_),
    .X(_0340_));
 sky130_fd_sc_hd__o21ai_2 _2368_ (.A1(_1337_),
    .A2(_0339_),
    .B1(_0340_),
    .Y(_0341_));
 sky130_fd_sc_hd__xnor2_1 _2369_ (.A(_0335_),
    .B(_0341_),
    .Y(_0342_));
 sky130_fd_sc_hd__xnor2_1 _2370_ (.A(_1337_),
    .B(_0339_),
    .Y(_0343_));
 sky130_fd_sc_hd__or2_1 _2371_ (.A(_0324_),
    .B(_0329_),
    .X(_0344_));
 sky130_fd_sc_hd__o21a_1 _2372_ (.A1(_1312_),
    .A2(_0330_),
    .B1(_0344_),
    .X(_0345_));
 sky130_fd_sc_hd__xnor2_2 _2373_ (.A(_0343_),
    .B(_0345_),
    .Y(_0346_));
 sky130_fd_sc_hd__or2_1 _2374_ (.A(_0342_),
    .B(_0346_),
    .X(_0347_));
 sky130_fd_sc_hd__nor2_1 _2375_ (.A(_0335_),
    .B(_0341_),
    .Y(_0348_));
 sky130_fd_sc_hd__or2_1 _2376_ (.A(_0343_),
    .B(_0345_),
    .X(_0349_));
 sky130_fd_sc_hd__or2b_1 _2377_ (.A(_0317_),
    .B_N(_0318_),
    .X(_0350_));
 sky130_fd_sc_hd__a21o_1 _2378_ (.A1(_0350_),
    .A2(_0333_),
    .B1(_0332_),
    .X(_0351_));
 sky130_fd_sc_hd__nand2_1 _2379_ (.A(_0335_),
    .B(_0341_),
    .Y(_0352_));
 sky130_fd_sc_hd__o221a_1 _2380_ (.A1(_0348_),
    .A2(_0349_),
    .B1(_0347_),
    .B2(_0351_),
    .C1(_0352_),
    .X(_0353_));
 sky130_fd_sc_hd__o31ai_4 _2381_ (.A1(_0320_),
    .A2(_0334_),
    .A3(_0347_),
    .B1(_0353_),
    .Y(_0354_));
 sky130_fd_sc_hd__xor2_2 _2382_ (.A(_1359_),
    .B(_1377_),
    .X(_0355_));
 sky130_fd_sc_hd__or2b_1 _2383_ (.A(_1412_),
    .B_N(_1414_),
    .X(_0356_));
 sky130_fd_sc_hd__xor2_2 _2384_ (.A(_0355_),
    .B(_0356_),
    .X(_0357_));
 sky130_fd_sc_hd__inv_2 _2385_ (.A(_1416_),
    .Y(_0358_));
 sky130_fd_sc_hd__a21oi_1 _2386_ (.A1(_0356_),
    .A2(_0358_),
    .B1(_0355_),
    .Y(_0359_));
 sky130_fd_sc_hd__a31o_1 _2387_ (.A1(_1418_),
    .A2(_0354_),
    .A3(_0357_),
    .B1(_0359_),
    .X(_0360_));
 sky130_fd_sc_hd__a21oi_2 _2388_ (.A1(_1382_),
    .A2(_0360_),
    .B1(_1380_),
    .Y(_0361_));
 sky130_fd_sc_hd__a31o_1 _2389_ (.A1(_1307_),
    .A2(net11),
    .A3(_1319_),
    .B1(_1318_),
    .X(_0362_));
 sky130_fd_sc_hd__xnor2_1 _2390_ (.A(_1408_),
    .B(_0362_),
    .Y(_0363_));
 sky130_fd_sc_hd__o21a_1 _2391_ (.A1(_1322_),
    .A2(_1325_),
    .B1(_0363_),
    .X(_0364_));
 sky130_fd_sc_hd__nor3_1 _2392_ (.A(_1322_),
    .B(_1325_),
    .C(_0363_),
    .Y(_0365_));
 sky130_fd_sc_hd__nor2_1 _2393_ (.A(_0364_),
    .B(_0365_),
    .Y(_0366_));
 sky130_fd_sc_hd__and2b_1 _2394_ (.A_N(_1343_),
    .B(_1327_),
    .X(_0367_));
 sky130_fd_sc_hd__and2_1 _2395_ (.A(_1309_),
    .B(_1344_),
    .X(_0368_));
 sky130_fd_sc_hd__nor2_1 _2396_ (.A(_0367_),
    .B(_0368_),
    .Y(_0369_));
 sky130_fd_sc_hd__xnor2_1 _2397_ (.A(_0366_),
    .B(_0369_),
    .Y(_0370_));
 sky130_fd_sc_hd__a21boi_2 _2398_ (.A1(_1357_),
    .A2(_0361_),
    .B1_N(_0370_),
    .Y(_0371_));
 sky130_fd_sc_hd__o21a_1 _2399_ (.A1(net14),
    .A2(_1320_),
    .B1(_1312_),
    .X(_0372_));
 sky130_fd_sc_hd__mux2_2 _2400_ (.A0(_1361_),
    .A1(_0372_),
    .S(_1338_),
    .X(_0373_));
 sky130_fd_sc_hd__o21ai_1 _2401_ (.A1(_0367_),
    .A2(_0368_),
    .B1(_0366_),
    .Y(_0374_));
 sky130_fd_sc_hd__and2b_1 _2402_ (.A_N(_0364_),
    .B(_0374_),
    .X(_0375_));
 sky130_fd_sc_hd__xnor2_2 _2403_ (.A(_0373_),
    .B(_0375_),
    .Y(_0376_));
 sky130_fd_sc_hd__o211a_1 _2404_ (.A1(_0367_),
    .A2(_0368_),
    .B1(_0366_),
    .C1(_0373_),
    .X(_0377_));
 sky130_fd_sc_hd__a21o_1 _2405_ (.A1(_0371_),
    .A2(_0376_),
    .B1(_0377_),
    .X(_0378_));
 sky130_fd_sc_hd__o21ai_1 _2406_ (.A1(net14),
    .A2(_1320_),
    .B1(_1319_),
    .Y(_0379_));
 sky130_fd_sc_hd__nand2_1 _2407_ (.A(_1338_),
    .B(_0379_),
    .Y(_0380_));
 sky130_fd_sc_hd__nand2_1 _2408_ (.A(_0364_),
    .B(_0373_),
    .Y(_0381_));
 sky130_fd_sc_hd__xor2_2 _2409_ (.A(_0380_),
    .B(_0381_),
    .X(_0382_));
 sky130_fd_sc_hd__nor2_1 _2410_ (.A(_1308_),
    .B(_1318_),
    .Y(_0383_));
 sky130_fd_sc_hd__nor2_1 _2411_ (.A(_0380_),
    .B(_0381_),
    .Y(_0384_));
 sky130_fd_sc_hd__a211oi_4 _2412_ (.A1(_0378_),
    .A2(_0382_),
    .B1(_0383_),
    .C1(_0384_),
    .Y(_0385_));
 sky130_fd_sc_hd__or2_1 _2413_ (.A(\simon0.play1.tick_counter[24] ),
    .B(_0385_),
    .X(_0386_));
 sky130_fd_sc_hd__inv_2 _2414_ (.A(\simon0.play1.tick_counter[23] ),
    .Y(_0387_));
 sky130_fd_sc_hd__xor2_2 _2415_ (.A(_0378_),
    .B(_0382_),
    .X(_0388_));
 sky130_fd_sc_hd__xor2_2 _2416_ (.A(_0371_),
    .B(_0376_),
    .X(_0389_));
 sky130_fd_sc_hd__inv_2 _2417_ (.A(\simon0.play1.tick_counter[22] ),
    .Y(_0390_));
 sky130_fd_sc_hd__a22oi_1 _2418_ (.A1(_0387_),
    .A2(_0388_),
    .B1(_0389_),
    .B2(_0390_),
    .Y(_0391_));
 sky130_fd_sc_hd__xnor2_2 _2419_ (.A(_1382_),
    .B(_0360_),
    .Y(_0392_));
 sky130_fd_sc_hd__inv_2 _2420_ (.A(\simon0.play1.tick_counter[21] ),
    .Y(_0393_));
 sky130_fd_sc_hd__xnor2_1 _2421_ (.A(_1357_),
    .B(_0370_),
    .Y(_0394_));
 sky130_fd_sc_hd__xnor2_2 _2422_ (.A(_0361_),
    .B(_0394_),
    .Y(_0395_));
 sky130_fd_sc_hd__a2bb2o_1 _2423_ (.A1_N(_0392_),
    .A2_N(\simon0.play1.tick_counter[20] ),
    .B1(_0393_),
    .B2(_0395_),
    .X(_0396_));
 sky130_fd_sc_hd__a211o_1 _2424_ (.A1(\simon0.play1.tick_counter[2] ),
    .A2(_0242_),
    .B1(\simon0.play1.tick_counter[0] ),
    .C1(\simon0.play1.tick_counter[1] ),
    .X(_0397_));
 sky130_fd_sc_hd__nand2_2 _2425_ (.A(_1307_),
    .B(net15),
    .Y(_0398_));
 sky130_fd_sc_hd__o22a_1 _2426_ (.A1(\simon0.play1.tick_counter[2] ),
    .A2(_0242_),
    .B1(_0398_),
    .B2(\simon0.play1.tick_counter[3] ),
    .X(_0399_));
 sky130_fd_sc_hd__xnor2_2 _2427_ (.A(_0290_),
    .B(_0296_),
    .Y(_0400_));
 sky130_fd_sc_hd__or3_1 _2428_ (.A(_0261_),
    .B(_0291_),
    .C(_0294_),
    .X(_0401_));
 sky130_fd_sc_hd__and2_1 _2429_ (.A(_0295_),
    .B(_0401_),
    .X(_0402_));
 sky130_fd_sc_hd__inv_2 _2430_ (.A(\simon0.play1.tick_counter[6] ),
    .Y(_0403_));
 sky130_fd_sc_hd__a2bb2o_1 _2431_ (.A1_N(\simon0.play1.tick_counter[7] ),
    .A2_N(_0400_),
    .B1(_0402_),
    .B2(_0403_),
    .X(_0404_));
 sky130_fd_sc_hd__nor2_1 _2432_ (.A(_0244_),
    .B(_0293_),
    .Y(_0405_));
 sky130_fd_sc_hd__or2_1 _2433_ (.A(_0294_),
    .B(_0405_),
    .X(_0406_));
 sky130_fd_sc_hd__a2bb2o_1 _2434_ (.A1_N(_0403_),
    .A2_N(_0402_),
    .B1(_0406_),
    .B2(\simon0.play1.tick_counter[5] ),
    .X(_0407_));
 sky130_fd_sc_hd__nand2_1 _2435_ (.A(\simon0.play1.tick_counter[7] ),
    .B(_0400_),
    .Y(_0408_));
 sky130_fd_sc_hd__or3b_1 _2436_ (.A(_0404_),
    .B(_0407_),
    .C_N(_0408_),
    .X(_0409_));
 sky130_fd_sc_hd__and2_1 _2437_ (.A(_0242_),
    .B(_0243_),
    .X(_0410_));
 sky130_fd_sc_hd__or2_1 _2438_ (.A(_0410_),
    .B(_0244_),
    .X(_0411_));
 sky130_fd_sc_hd__and2_1 _2439_ (.A(\simon0.play1.tick_counter[4] ),
    .B(_0411_),
    .X(_0412_));
 sky130_fd_sc_hd__o22a_1 _2440_ (.A1(\simon0.play1.tick_counter[5] ),
    .A2(_0406_),
    .B1(_0411_),
    .B2(\simon0.play1.tick_counter[4] ),
    .X(_0413_));
 sky130_fd_sc_hd__or3b_1 _2441_ (.A(_0409_),
    .B(_0412_),
    .C_N(_0413_),
    .X(_0414_));
 sky130_fd_sc_hd__and2_1 _2442_ (.A(\simon0.play1.tick_counter[3] ),
    .B(_0398_),
    .X(_0415_));
 sky130_fd_sc_hd__a211o_1 _2443_ (.A1(_0397_),
    .A2(_0399_),
    .B1(_0414_),
    .C1(_0415_),
    .X(_0416_));
 sky130_fd_sc_hd__o2bb2a_1 _2444_ (.A1_N(_0408_),
    .A2_N(_0404_),
    .B1(_0409_),
    .B2(_0413_),
    .X(_0417_));
 sky130_fd_sc_hd__nor2b_1 _2445_ (.A(_0271_),
    .B_N(_0270_),
    .Y(_0418_));
 sky130_fd_sc_hd__and2_1 _2446_ (.A(_0267_),
    .B(_0302_),
    .X(_0419_));
 sky130_fd_sc_hd__a21bo_1 _2447_ (.A1(_0301_),
    .A2(_0419_),
    .B1_N(_0267_),
    .X(_0420_));
 sky130_fd_sc_hd__xnor2_1 _2448_ (.A(_0418_),
    .B(_0420_),
    .Y(_0421_));
 sky130_fd_sc_hd__xnor2_2 _2449_ (.A(_0301_),
    .B(_0419_),
    .Y(_0422_));
 sky130_fd_sc_hd__o22a_1 _2450_ (.A1(\simon0.play1.tick_counter[11] ),
    .A2(_0421_),
    .B1(_0422_),
    .B2(\simon0.play1.tick_counter[10] ),
    .X(_0423_));
 sky130_fd_sc_hd__nand2_1 _2451_ (.A(\simon0.play1.tick_counter[10] ),
    .B(_0422_),
    .Y(_0424_));
 sky130_fd_sc_hd__nand2_1 _2452_ (.A(\simon0.play1.tick_counter[11] ),
    .B(_0421_),
    .Y(_0425_));
 sky130_fd_sc_hd__nand3_1 _2453_ (.A(_0423_),
    .B(_0424_),
    .C(_0425_),
    .Y(_0426_));
 sky130_fd_sc_hd__xnor2_2 _2454_ (.A(_0289_),
    .B(_0297_),
    .Y(_0427_));
 sky130_fd_sc_hd__and2_1 _2455_ (.A(\simon0.play1.tick_counter[8] ),
    .B(_0427_),
    .X(_0428_));
 sky130_fd_sc_hd__and3_1 _2456_ (.A(_0300_),
    .B(_0285_),
    .C(_0299_),
    .X(_0429_));
 sky130_fd_sc_hd__a21oi_1 _2457_ (.A1(_0300_),
    .A2(_0285_),
    .B1(_0299_),
    .Y(_0430_));
 sky130_fd_sc_hd__or2_1 _2458_ (.A(_0429_),
    .B(_0430_),
    .X(_0431_));
 sky130_fd_sc_hd__and2_1 _2459_ (.A(\simon0.play1.tick_counter[9] ),
    .B(_0431_),
    .X(_0432_));
 sky130_fd_sc_hd__o22a_1 _2460_ (.A1(\simon0.play1.tick_counter[8] ),
    .A2(_0427_),
    .B1(_0431_),
    .B2(\simon0.play1.tick_counter[9] ),
    .X(_0433_));
 sky130_fd_sc_hd__or4b_1 _2461_ (.A(_0426_),
    .B(_0428_),
    .C(_0432_),
    .D_N(_0433_),
    .X(_0434_));
 sky130_fd_sc_hd__inv_2 _2462_ (.A(\simon0.play1.tick_counter[15] ),
    .Y(_0435_));
 sky130_fd_sc_hd__a21o_1 _2463_ (.A1(_0350_),
    .A2(_0320_),
    .B1(_0334_),
    .X(_0436_));
 sky130_fd_sc_hd__nand3_1 _2464_ (.A(_0350_),
    .B(_0320_),
    .C(_0334_),
    .Y(_0437_));
 sky130_fd_sc_hd__nand4_1 _2465_ (.A(_0319_),
    .B(_0233_),
    .C(_0274_),
    .D(_0304_),
    .Y(_0438_));
 sky130_fd_sc_hd__and2_1 _2466_ (.A(_0320_),
    .B(_0438_),
    .X(_0439_));
 sky130_fd_sc_hd__inv_2 _2467_ (.A(\simon0.play1.tick_counter[14] ),
    .Y(_0440_));
 sky130_fd_sc_hd__a32o_1 _2468_ (.A1(_0435_),
    .A2(_0436_),
    .A3(_0437_),
    .B1(_0439_),
    .B2(_0440_),
    .X(_0441_));
 sky130_fd_sc_hd__a21o_1 _2469_ (.A1(_0301_),
    .A2(_0303_),
    .B1(_0272_),
    .X(_0442_));
 sky130_fd_sc_hd__xnor2_2 _2470_ (.A(_0234_),
    .B(_0442_),
    .Y(_0443_));
 sky130_fd_sc_hd__inv_2 _2471_ (.A(\simon0.play1.tick_counter[13] ),
    .Y(_0444_));
 sky130_fd_sc_hd__a21boi_1 _2472_ (.A1(_0234_),
    .A2(_0442_),
    .B1_N(_0231_),
    .Y(_0445_));
 sky130_fd_sc_hd__xnor2_1 _2473_ (.A(_0445_),
    .B(_0273_),
    .Y(_0446_));
 sky130_fd_sc_hd__a2bb2o_1 _2474_ (.A1_N(_0443_),
    .A2_N(\simon0.play1.tick_counter[12] ),
    .B1(_0444_),
    .B2(_0446_),
    .X(_0447_));
 sky130_fd_sc_hd__a21o_1 _2475_ (.A1(_0436_),
    .A2(_0437_),
    .B1(_0435_),
    .X(_0448_));
 sky130_fd_sc_hd__nand2_1 _2476_ (.A(\simon0.play1.tick_counter[12] ),
    .B(_0443_),
    .Y(_0449_));
 sky130_fd_sc_hd__o221a_1 _2477_ (.A1(_0440_),
    .A2(_0439_),
    .B1(_0446_),
    .B2(_0444_),
    .C1(_0449_),
    .X(_0450_));
 sky130_fd_sc_hd__or4bb_2 _2478_ (.A(_0441_),
    .B(_0447_),
    .C_N(_0448_),
    .D_N(_0450_),
    .X(_0451_));
 sky130_fd_sc_hd__a211oi_2 _2479_ (.A1(_0416_),
    .A2(_0417_),
    .B1(_0434_),
    .C1(_0451_),
    .Y(_0452_));
 sky130_fd_sc_hd__inv_2 _2480_ (.A(_0425_),
    .Y(_0453_));
 sky130_fd_sc_hd__o32a_1 _2481_ (.A1(_0426_),
    .A2(_0433_),
    .A3(_0432_),
    .B1(_0453_),
    .B2(_0423_),
    .X(_0454_));
 sky130_fd_sc_hd__o22a_1 _2482_ (.A1(_0440_),
    .A2(_0439_),
    .B1(_0446_),
    .B2(_0444_),
    .X(_0455_));
 sky130_fd_sc_hd__a21o_1 _2483_ (.A1(_0455_),
    .A2(_0447_),
    .B1(_0441_),
    .X(_0456_));
 sky130_fd_sc_hd__a2bb2o_1 _2484_ (.A1_N(_0451_),
    .A2_N(_0454_),
    .B1(_0456_),
    .B2(_0448_),
    .X(_0457_));
 sky130_fd_sc_hd__inv_2 _2485_ (.A(\simon0.play1.tick_counter[19] ),
    .Y(_0458_));
 sky130_fd_sc_hd__a21oi_1 _2486_ (.A1(_1418_),
    .A2(_0354_),
    .B1(_1416_),
    .Y(_0459_));
 sky130_fd_sc_hd__xnor2_2 _2487_ (.A(_0357_),
    .B(_0459_),
    .Y(_0460_));
 sky130_fd_sc_hd__o21ai_1 _2488_ (.A1(_0320_),
    .A2(_0334_),
    .B1(_0351_),
    .Y(_0461_));
 sky130_fd_sc_hd__xor2_2 _2489_ (.A(_0346_),
    .B(_0461_),
    .X(_0462_));
 sky130_fd_sc_hd__nand2_1 _2490_ (.A(\simon0.play1.tick_counter[16] ),
    .B(_0462_),
    .Y(_0463_));
 sky130_fd_sc_hd__a311o_1 _2491_ (.A1(_0350_),
    .A2(_0320_),
    .A3(_0333_),
    .B1(_0346_),
    .C1(_0332_),
    .X(_0464_));
 sky130_fd_sc_hd__nand3b_1 _2492_ (.A_N(_0342_),
    .B(_0349_),
    .C(_0464_),
    .Y(_0465_));
 sky130_fd_sc_hd__a21bo_1 _2493_ (.A1(_0349_),
    .A2(_0464_),
    .B1_N(_0342_),
    .X(_0466_));
 sky130_fd_sc_hd__xnor2_2 _2494_ (.A(_1418_),
    .B(_0354_),
    .Y(_0467_));
 sky130_fd_sc_hd__a32oi_1 _2495_ (.A1(\simon0.play1.tick_counter[17] ),
    .A2(_0465_),
    .A3(_0466_),
    .B1(_0467_),
    .B2(\simon0.play1.tick_counter[18] ),
    .Y(_0468_));
 sky130_fd_sc_hd__o211a_1 _2496_ (.A1(_0458_),
    .A2(_0460_),
    .B1(_0463_),
    .C1(_0468_),
    .X(_0469_));
 sky130_fd_sc_hd__a21oi_1 _2497_ (.A1(_0349_),
    .A2(_0464_),
    .B1(_0342_),
    .Y(_0470_));
 sky130_fd_sc_hd__and3_1 _2498_ (.A(_0342_),
    .B(_0349_),
    .C(_0464_),
    .X(_0471_));
 sky130_fd_sc_hd__o32a_1 _2499_ (.A1(\simon0.play1.tick_counter[17] ),
    .A2(_0470_),
    .A3(_0471_),
    .B1(_0462_),
    .B2(\simon0.play1.tick_counter[16] ),
    .X(_0472_));
 sky130_fd_sc_hd__o2bb2a_1 _2500_ (.A1_N(_0458_),
    .A2_N(_0460_),
    .B1(_0467_),
    .B2(\simon0.play1.tick_counter[18] ),
    .X(_0473_));
 sky130_fd_sc_hd__o2111a_1 _2501_ (.A1(_0452_),
    .A2(_0457_),
    .B1(_0469_),
    .C1(_0472_),
    .D1(_0473_),
    .X(_0474_));
 sky130_fd_sc_hd__or2b_1 _2502_ (.A(_0472_),
    .B_N(_0468_),
    .X(_0475_));
 sky130_fd_sc_hd__o2bb2a_1 _2503_ (.A1_N(_0473_),
    .A2_N(_0475_),
    .B1(_0458_),
    .B2(_0460_),
    .X(_0476_));
 sky130_fd_sc_hd__nand2_1 _2504_ (.A(\simon0.play1.tick_counter[20] ),
    .B(_0392_),
    .Y(_0477_));
 sky130_fd_sc_hd__or3b_1 _2505_ (.A(_0397_),
    .B(_0415_),
    .C_N(_0399_),
    .X(_0478_));
 sky130_fd_sc_hd__nor4_1 _2506_ (.A(_0434_),
    .B(_0451_),
    .C(_0414_),
    .D(_0478_),
    .Y(_0479_));
 sky130_fd_sc_hd__nand4_1 _2507_ (.A(_0469_),
    .B(_0472_),
    .C(_0473_),
    .D(_0479_),
    .Y(_0480_));
 sky130_fd_sc_hd__o211a_1 _2508_ (.A1(_0474_),
    .A2(_0476_),
    .B1(_0477_),
    .C1(_0480_),
    .X(_0481_));
 sky130_fd_sc_hd__o22a_1 _2509_ (.A1(_0390_),
    .A2(_0389_),
    .B1(_0395_),
    .B2(_0393_),
    .X(_0482_));
 sky130_fd_sc_hd__o21ai_1 _2510_ (.A1(_0396_),
    .A2(_0481_),
    .B1(_0482_),
    .Y(_0483_));
 sky130_fd_sc_hd__nor2_1 _2511_ (.A(_0387_),
    .B(_0388_),
    .Y(_0484_));
 sky130_fd_sc_hd__a221o_1 _2512_ (.A1(\simon0.play1.tick_counter[24] ),
    .A2(_0385_),
    .B1(_0391_),
    .B2(_0483_),
    .C1(_0484_),
    .X(_0485_));
 sky130_fd_sc_hd__or4_1 _2513_ (.A(\simon0.play1.tick_counter[31] ),
    .B(\simon0.play1.tick_counter[30] ),
    .C(\simon0.play1.tick_counter[29] ),
    .D(\simon0.play1.tick_counter[28] ),
    .X(_0486_));
 sky130_fd_sc_hd__or4_2 _2514_ (.A(\simon0.play1.tick_counter[27] ),
    .B(\simon0.play1.tick_counter[26] ),
    .C(\simon0.play1.tick_counter[25] ),
    .D(_0486_),
    .X(_0487_));
 sky130_fd_sc_hd__a21oi_4 _2515_ (.A1(_0386_),
    .A2(_0485_),
    .B1(_0487_),
    .Y(_0488_));
 sky130_fd_sc_hd__clkbuf_4 _2516_ (.A(_0488_),
    .X(_0489_));
 sky130_fd_sc_hd__nor2_2 _2517_ (.A(\simon0.play1.freq[2] ),
    .B(\simon0.play1.tick_counter[2] ),
    .Y(_0490_));
 sky130_fd_sc_hd__and2_1 _2518_ (.A(\simon0.play1.freq[2] ),
    .B(\simon0.play1.tick_counter[2] ),
    .X(_0491_));
 sky130_fd_sc_hd__nor2_1 _2519_ (.A(_0490_),
    .B(_0491_),
    .Y(_0492_));
 sky130_fd_sc_hd__and2_1 _2520_ (.A(\simon0.play1.freq[1] ),
    .B(\simon0.play1.tick_counter[1] ),
    .X(_0493_));
 sky130_fd_sc_hd__a21oi_1 _2521_ (.A1(_1295_),
    .A2(_1296_),
    .B1(_0493_),
    .Y(_0494_));
 sky130_fd_sc_hd__xnor2_1 _2522_ (.A(_0492_),
    .B(_0494_),
    .Y(_0495_));
 sky130_fd_sc_hd__or2_1 _2523_ (.A(_0242_),
    .B(_0495_),
    .X(_0496_));
 sky130_fd_sc_hd__o21ai_1 _2524_ (.A1(_0489_),
    .A2(_0496_),
    .B1(_1302_),
    .Y(_0497_));
 sky130_fd_sc_hd__o21a_1 _2525_ (.A1(_0242_),
    .A2(_0488_),
    .B1(_0495_),
    .X(_0498_));
 sky130_fd_sc_hd__clkbuf_4 _2526_ (.A(_1084_),
    .X(_0499_));
 sky130_fd_sc_hd__o221a_1 _2527_ (.A1(\simon0.play1.tick_counter[2] ),
    .A2(_1303_),
    .B1(_0497_),
    .B2(_0498_),
    .C1(_0499_),
    .X(_0049_));
 sky130_fd_sc_hd__a21o_1 _2528_ (.A1(_0386_),
    .A2(_0485_),
    .B1(_0487_),
    .X(_0500_));
 sky130_fd_sc_hd__clkbuf_4 _2529_ (.A(_0500_),
    .X(_0501_));
 sky130_fd_sc_hd__clkbuf_4 _2530_ (.A(_0501_),
    .X(_0502_));
 sky130_fd_sc_hd__nor2_1 _2531_ (.A(\simon0.play1.freq[3] ),
    .B(\simon0.play1.tick_counter[3] ),
    .Y(_0503_));
 sky130_fd_sc_hd__nand2_1 _2532_ (.A(\simon0.play1.freq[3] ),
    .B(\simon0.play1.tick_counter[3] ),
    .Y(_0504_));
 sky130_fd_sc_hd__or2b_1 _2533_ (.A(_0503_),
    .B_N(_0504_),
    .X(_0505_));
 sky130_fd_sc_hd__a211oi_4 _2534_ (.A1(_1295_),
    .A2(_1296_),
    .B1(_0491_),
    .C1(_0493_),
    .Y(_0506_));
 sky130_fd_sc_hd__or2_1 _2535_ (.A(_0490_),
    .B(_0506_),
    .X(_0507_));
 sky130_fd_sc_hd__xnor2_2 _2536_ (.A(_0505_),
    .B(_0507_),
    .Y(_0508_));
 sky130_fd_sc_hd__nor2_1 _2537_ (.A(_0502_),
    .B(_0508_),
    .Y(_0509_));
 sky130_fd_sc_hd__clkbuf_4 _2538_ (.A(_0501_),
    .X(_0510_));
 sky130_fd_sc_hd__xnor2_1 _2539_ (.A(_0398_),
    .B(_0508_),
    .Y(_0511_));
 sky130_fd_sc_hd__nand2_1 _2540_ (.A(_0496_),
    .B(_0511_),
    .Y(_0512_));
 sky130_fd_sc_hd__or2_1 _2541_ (.A(_0496_),
    .B(_0511_),
    .X(_0513_));
 sky130_fd_sc_hd__nor4_4 _2542_ (.A(\simon0.play1.freq[9] ),
    .B(\simon0.play1.freq[8] ),
    .C(_1298_),
    .D(_1299_),
    .Y(_0514_));
 sky130_fd_sc_hd__a31o_1 _2543_ (.A1(_0510_),
    .A2(_0512_),
    .A3(_0513_),
    .B1(_0514_),
    .X(_0515_));
 sky130_fd_sc_hd__o221a_1 _2544_ (.A1(\simon0.play1.tick_counter[3] ),
    .A2(_1303_),
    .B1(_0509_),
    .B2(_0515_),
    .C1(_0499_),
    .X(_0050_));
 sky130_fd_sc_hd__or2_1 _2545_ (.A(\simon0.play1.freq[4] ),
    .B(\simon0.play1.tick_counter[4] ),
    .X(_0516_));
 sky130_fd_sc_hd__nand2_1 _2546_ (.A(\simon0.play1.freq[4] ),
    .B(\simon0.play1.tick_counter[4] ),
    .Y(_0517_));
 sky130_fd_sc_hd__nand2_1 _2547_ (.A(_0516_),
    .B(_0517_),
    .Y(_0518_));
 sky130_fd_sc_hd__o31a_1 _2548_ (.A1(_0490_),
    .A2(_0503_),
    .A3(_0506_),
    .B1(_0504_),
    .X(_0519_));
 sky130_fd_sc_hd__xnor2_1 _2549_ (.A(_0518_),
    .B(_0519_),
    .Y(_0520_));
 sky130_fd_sc_hd__nor2_1 _2550_ (.A(_0502_),
    .B(_0520_),
    .Y(_0521_));
 sky130_fd_sc_hd__nor2_1 _2551_ (.A(_0410_),
    .B(_0244_),
    .Y(_0522_));
 sky130_fd_sc_hd__nand2_1 _2552_ (.A(_0522_),
    .B(_0520_),
    .Y(_0523_));
 sky130_fd_sc_hd__or2_1 _2553_ (.A(_0522_),
    .B(_0520_),
    .X(_0524_));
 sky130_fd_sc_hd__nand2_1 _2554_ (.A(_0523_),
    .B(_0524_),
    .Y(_0525_));
 sky130_fd_sc_hd__a21oi_1 _2555_ (.A1(_1307_),
    .A2(net15),
    .B1(_0508_),
    .Y(_0526_));
 sky130_fd_sc_hd__a21o_1 _2556_ (.A1(_0496_),
    .A2(_0511_),
    .B1(_0526_),
    .X(_0527_));
 sky130_fd_sc_hd__xnor2_1 _2557_ (.A(_0525_),
    .B(_0527_),
    .Y(_0528_));
 sky130_fd_sc_hd__clkbuf_4 _2558_ (.A(_0514_),
    .X(_0529_));
 sky130_fd_sc_hd__a21o_1 _2559_ (.A1(_0510_),
    .A2(_0528_),
    .B1(_0529_),
    .X(_0530_));
 sky130_fd_sc_hd__o221a_1 _2560_ (.A1(\simon0.play1.tick_counter[4] ),
    .A2(_1303_),
    .B1(_0521_),
    .B2(_0530_),
    .C1(_0499_),
    .X(_0051_));
 sky130_fd_sc_hd__or2_1 _2561_ (.A(\simon0.play1.freq[5] ),
    .B(\simon0.play1.tick_counter[5] ),
    .X(_0531_));
 sky130_fd_sc_hd__nand2_1 _2562_ (.A(\simon0.play1.freq[5] ),
    .B(\simon0.play1.tick_counter[5] ),
    .Y(_0532_));
 sky130_fd_sc_hd__nand2_1 _2563_ (.A(_0531_),
    .B(_0532_),
    .Y(_0533_));
 sky130_fd_sc_hd__o311ai_4 _2564_ (.A1(_0490_),
    .A2(_0503_),
    .A3(_0506_),
    .B1(_0517_),
    .C1(_0504_),
    .Y(_0534_));
 sky130_fd_sc_hd__nand2_1 _2565_ (.A(_0516_),
    .B(_0534_),
    .Y(_0535_));
 sky130_fd_sc_hd__xor2_1 _2566_ (.A(_0533_),
    .B(_0535_),
    .X(_0536_));
 sky130_fd_sc_hd__nor2_1 _2567_ (.A(_0406_),
    .B(_0536_),
    .Y(_0537_));
 sky130_fd_sc_hd__nand2_1 _2568_ (.A(_0406_),
    .B(_0536_),
    .Y(_0538_));
 sky130_fd_sc_hd__or2b_1 _2569_ (.A(_0537_),
    .B_N(_0538_),
    .X(_0539_));
 sky130_fd_sc_hd__nand2_1 _2570_ (.A(_0523_),
    .B(_0527_),
    .Y(_0540_));
 sky130_fd_sc_hd__nand2_1 _2571_ (.A(_0524_),
    .B(_0540_),
    .Y(_0541_));
 sky130_fd_sc_hd__xnor2_1 _2572_ (.A(_0539_),
    .B(_0541_),
    .Y(_0542_));
 sky130_fd_sc_hd__mux2_1 _2573_ (.A0(_0536_),
    .A1(_0542_),
    .S(_0501_),
    .X(_0543_));
 sky130_fd_sc_hd__or2_1 _2574_ (.A(\simon0.play1.tick_counter[5] ),
    .B(_1302_),
    .X(_0544_));
 sky130_fd_sc_hd__o211a_1 _2575_ (.A1(_0529_),
    .A2(_0543_),
    .B1(_0544_),
    .C1(_1190_),
    .X(_0052_));
 sky130_fd_sc_hd__nor2_1 _2576_ (.A(\simon0.play1.freq[6] ),
    .B(\simon0.play1.tick_counter[6] ),
    .Y(_0545_));
 sky130_fd_sc_hd__nand2_1 _2577_ (.A(\simon0.play1.freq[6] ),
    .B(\simon0.play1.tick_counter[6] ),
    .Y(_0546_));
 sky130_fd_sc_hd__or2b_1 _2578_ (.A(_0545_),
    .B_N(_0546_),
    .X(_0547_));
 sky130_fd_sc_hd__and2_1 _2579_ (.A(\simon0.play1.freq[5] ),
    .B(\simon0.play1.tick_counter[5] ),
    .X(_0548_));
 sky130_fd_sc_hd__a31oi_2 _2580_ (.A1(_0516_),
    .A2(_0531_),
    .A3(_0534_),
    .B1(_0548_),
    .Y(_0549_));
 sky130_fd_sc_hd__xnor2_1 _2581_ (.A(_0547_),
    .B(_0549_),
    .Y(_0550_));
 sky130_fd_sc_hd__nor2_1 _2582_ (.A(_0502_),
    .B(_0550_),
    .Y(_0551_));
 sky130_fd_sc_hd__nand2_1 _2583_ (.A(_0402_),
    .B(_0550_),
    .Y(_0552_));
 sky130_fd_sc_hd__or2_1 _2584_ (.A(_0402_),
    .B(_0550_),
    .X(_0553_));
 sky130_fd_sc_hd__nand2_1 _2585_ (.A(_0552_),
    .B(_0553_),
    .Y(_0554_));
 sky130_fd_sc_hd__a31o_1 _2586_ (.A1(_0524_),
    .A2(_0538_),
    .A3(_0540_),
    .B1(_0537_),
    .X(_0555_));
 sky130_fd_sc_hd__xor2_1 _2587_ (.A(_0554_),
    .B(_0555_),
    .X(_0556_));
 sky130_fd_sc_hd__a21o_1 _2588_ (.A1(_0510_),
    .A2(_0556_),
    .B1(_0529_),
    .X(_0557_));
 sky130_fd_sc_hd__o221a_1 _2589_ (.A1(\simon0.play1.tick_counter[6] ),
    .A2(_1303_),
    .B1(_0551_),
    .B2(_0557_),
    .C1(_0499_),
    .X(_0053_));
 sky130_fd_sc_hd__or2_1 _2590_ (.A(\simon0.play1.freq[7] ),
    .B(\simon0.play1.tick_counter[7] ),
    .X(_0558_));
 sky130_fd_sc_hd__nand2_1 _2591_ (.A(\simon0.play1.freq[7] ),
    .B(\simon0.play1.tick_counter[7] ),
    .Y(_0559_));
 sky130_fd_sc_hd__nand2_1 _2592_ (.A(_0558_),
    .B(_0559_),
    .Y(_0560_));
 sky130_fd_sc_hd__o21ai_2 _2593_ (.A1(_0545_),
    .A2(_0549_),
    .B1(_0546_),
    .Y(_0561_));
 sky130_fd_sc_hd__xnor2_1 _2594_ (.A(_0560_),
    .B(_0561_),
    .Y(_0562_));
 sky130_fd_sc_hd__or2_1 _2595_ (.A(_0400_),
    .B(_0562_),
    .X(_0563_));
 sky130_fd_sc_hd__nand2_1 _2596_ (.A(_0400_),
    .B(_0562_),
    .Y(_0564_));
 sky130_fd_sc_hd__nand2_1 _2597_ (.A(_0563_),
    .B(_0564_),
    .Y(_0565_));
 sky130_fd_sc_hd__o21a_1 _2598_ (.A1(_0554_),
    .A2(_0555_),
    .B1(_0553_),
    .X(_0566_));
 sky130_fd_sc_hd__xnor2_1 _2599_ (.A(_0565_),
    .B(_0566_),
    .Y(_0567_));
 sky130_fd_sc_hd__nor2_1 _2600_ (.A(_0489_),
    .B(_0567_),
    .Y(_0568_));
 sky130_fd_sc_hd__a21o_1 _2601_ (.A1(_0489_),
    .A2(_0562_),
    .B1(_0529_),
    .X(_0569_));
 sky130_fd_sc_hd__o221a_1 _2602_ (.A1(\simon0.play1.tick_counter[7] ),
    .A2(_1303_),
    .B1(_0568_),
    .B2(_0569_),
    .C1(_0499_),
    .X(_0054_));
 sky130_fd_sc_hd__clkbuf_4 _2603_ (.A(_1302_),
    .X(_0570_));
 sky130_fd_sc_hd__nor2_1 _2604_ (.A(\simon0.play1.freq[8] ),
    .B(\simon0.play1.tick_counter[8] ),
    .Y(_0571_));
 sky130_fd_sc_hd__nand2_1 _2605_ (.A(\simon0.play1.freq[8] ),
    .B(\simon0.play1.tick_counter[8] ),
    .Y(_0572_));
 sky130_fd_sc_hd__or2b_1 _2606_ (.A(_0571_),
    .B_N(_0572_),
    .X(_0573_));
 sky130_fd_sc_hd__a21boi_4 _2607_ (.A1(_0558_),
    .A2(_0561_),
    .B1_N(_0559_),
    .Y(_0574_));
 sky130_fd_sc_hd__xor2_2 _2608_ (.A(_0573_),
    .B(_0574_),
    .X(_0575_));
 sky130_fd_sc_hd__xnor2_1 _2609_ (.A(_0427_),
    .B(_0575_),
    .Y(_0576_));
 sky130_fd_sc_hd__o211ai_1 _2610_ (.A1(_0554_),
    .A2(_0555_),
    .B1(_0564_),
    .C1(_0553_),
    .Y(_0577_));
 sky130_fd_sc_hd__nand2_1 _2611_ (.A(_0563_),
    .B(_0577_),
    .Y(_0578_));
 sky130_fd_sc_hd__xnor2_1 _2612_ (.A(_0576_),
    .B(_0578_),
    .Y(_0579_));
 sky130_fd_sc_hd__nor2_1 _2613_ (.A(_0489_),
    .B(_0579_),
    .Y(_0580_));
 sky130_fd_sc_hd__a21o_1 _2614_ (.A1(_0489_),
    .A2(_0575_),
    .B1(_0529_),
    .X(_0581_));
 sky130_fd_sc_hd__o221a_1 _2615_ (.A1(\simon0.play1.tick_counter[8] ),
    .A2(_0570_),
    .B1(_0580_),
    .B2(_0581_),
    .C1(_0499_),
    .X(_0055_));
 sky130_fd_sc_hd__or2_1 _2616_ (.A(\simon0.play1.freq[9] ),
    .B(\simon0.play1.tick_counter[9] ),
    .X(_0582_));
 sky130_fd_sc_hd__nand2_1 _2617_ (.A(\simon0.play1.freq[9] ),
    .B(\simon0.play1.tick_counter[9] ),
    .Y(_0583_));
 sky130_fd_sc_hd__nand2_1 _2618_ (.A(_0582_),
    .B(_0583_),
    .Y(_0584_));
 sky130_fd_sc_hd__o21ai_1 _2619_ (.A1(_0571_),
    .A2(_0574_),
    .B1(_0572_),
    .Y(_0585_));
 sky130_fd_sc_hd__xnor2_1 _2620_ (.A(_0584_),
    .B(_0585_),
    .Y(_0586_));
 sky130_fd_sc_hd__nor2_1 _2621_ (.A(_0431_),
    .B(_0586_),
    .Y(_0587_));
 sky130_fd_sc_hd__o21a_1 _2622_ (.A1(_0429_),
    .A2(_0430_),
    .B1(_0586_),
    .X(_0588_));
 sky130_fd_sc_hd__or2_1 _2623_ (.A(_0587_),
    .B(_0588_),
    .X(_0589_));
 sky130_fd_sc_hd__a22o_1 _2624_ (.A1(_0427_),
    .A2(_0575_),
    .B1(_0577_),
    .B2(_0563_),
    .X(_0590_));
 sky130_fd_sc_hd__o21a_1 _2625_ (.A1(_0427_),
    .A2(_0575_),
    .B1(_0590_),
    .X(_0591_));
 sky130_fd_sc_hd__xnor2_1 _2626_ (.A(_0589_),
    .B(_0591_),
    .Y(_0592_));
 sky130_fd_sc_hd__mux2_1 _2627_ (.A0(_0586_),
    .A1(_0592_),
    .S(_0501_),
    .X(_0593_));
 sky130_fd_sc_hd__or2_1 _2628_ (.A(\simon0.play1.tick_counter[9] ),
    .B(_1302_),
    .X(_0594_));
 sky130_fd_sc_hd__o211a_1 _2629_ (.A1(_0529_),
    .A2(_0593_),
    .B1(_0594_),
    .C1(_1190_),
    .X(_0056_));
 sky130_fd_sc_hd__clkbuf_4 _2630_ (.A(_1301_),
    .X(_0595_));
 sky130_fd_sc_hd__o211ai_2 _2631_ (.A1(_0571_),
    .A2(_0574_),
    .B1(_0583_),
    .C1(_0572_),
    .Y(_0596_));
 sky130_fd_sc_hd__nand2_1 _2632_ (.A(_0582_),
    .B(_0596_),
    .Y(_0597_));
 sky130_fd_sc_hd__xor2_1 _2633_ (.A(\simon0.play1.tick_counter[10] ),
    .B(_0597_),
    .X(_0598_));
 sky130_fd_sc_hd__xnor2_1 _2634_ (.A(_0422_),
    .B(_0598_),
    .Y(_0599_));
 sky130_fd_sc_hd__o32a_1 _2635_ (.A1(_0429_),
    .A2(_0430_),
    .A3(_0586_),
    .B1(_0588_),
    .B2(_0591_),
    .X(_0600_));
 sky130_fd_sc_hd__and2_1 _2636_ (.A(_0599_),
    .B(_0600_),
    .X(_0601_));
 sky130_fd_sc_hd__nor2_1 _2637_ (.A(_0599_),
    .B(_0600_),
    .Y(_0602_));
 sky130_fd_sc_hd__or2_1 _2638_ (.A(_0501_),
    .B(_0598_),
    .X(_0603_));
 sky130_fd_sc_hd__o31a_1 _2639_ (.A1(_0488_),
    .A2(_0601_),
    .A3(_0602_),
    .B1(_0603_),
    .X(_0604_));
 sky130_fd_sc_hd__nand2_1 _2640_ (.A(_0595_),
    .B(_0604_),
    .Y(_0605_));
 sky130_fd_sc_hd__o211a_1 _2641_ (.A1(\simon0.play1.tick_counter[10] ),
    .A2(_1303_),
    .B1(_0605_),
    .C1(_1190_),
    .X(_0057_));
 sky130_fd_sc_hd__and4_1 _2642_ (.A(\simon0.play1.tick_counter[11] ),
    .B(\simon0.play1.tick_counter[10] ),
    .C(_0582_),
    .D(_0596_),
    .X(_0606_));
 sky130_fd_sc_hd__a31o_1 _2643_ (.A1(\simon0.play1.tick_counter[10] ),
    .A2(_0582_),
    .A3(_0596_),
    .B1(\simon0.play1.tick_counter[11] ),
    .X(_0607_));
 sky130_fd_sc_hd__nand2b_1 _2644_ (.A_N(_0606_),
    .B(_0607_),
    .Y(_0608_));
 sky130_fd_sc_hd__nor2_1 _2645_ (.A(_0502_),
    .B(_0608_),
    .Y(_0609_));
 sky130_fd_sc_hd__and2b_1 _2646_ (.A_N(_0598_),
    .B(_0422_),
    .X(_0610_));
 sky130_fd_sc_hd__nor2_1 _2647_ (.A(_0610_),
    .B(_0601_),
    .Y(_0611_));
 sky130_fd_sc_hd__xor2_1 _2648_ (.A(_0418_),
    .B(_0420_),
    .X(_0612_));
 sky130_fd_sc_hd__nor2_1 _2649_ (.A(_0612_),
    .B(_0608_),
    .Y(_0613_));
 sky130_fd_sc_hd__nand2_1 _2650_ (.A(_0612_),
    .B(_0608_),
    .Y(_0614_));
 sky130_fd_sc_hd__or2b_1 _2651_ (.A(_0613_),
    .B_N(_0614_),
    .X(_0615_));
 sky130_fd_sc_hd__xnor2_1 _2652_ (.A(_0611_),
    .B(_0615_),
    .Y(_0616_));
 sky130_fd_sc_hd__o21ai_1 _2653_ (.A1(_0489_),
    .A2(_0616_),
    .B1(_1302_),
    .Y(_0617_));
 sky130_fd_sc_hd__clkbuf_4 _2654_ (.A(_1084_),
    .X(_0618_));
 sky130_fd_sc_hd__o221a_1 _2655_ (.A1(\simon0.play1.tick_counter[11] ),
    .A2(_0570_),
    .B1(_0609_),
    .B2(_0617_),
    .C1(_0618_),
    .X(_0058_));
 sky130_fd_sc_hd__xnor2_1 _2656_ (.A(\simon0.play1.tick_counter[12] ),
    .B(_0606_),
    .Y(_0619_));
 sky130_fd_sc_hd__nor2_1 _2657_ (.A(_0502_),
    .B(_0619_),
    .Y(_0620_));
 sky130_fd_sc_hd__o21a_1 _2658_ (.A1(_0610_),
    .A2(_0601_),
    .B1(_0614_),
    .X(_0621_));
 sky130_fd_sc_hd__xnor2_1 _2659_ (.A(_0443_),
    .B(_0619_),
    .Y(_0622_));
 sky130_fd_sc_hd__o21ai_1 _2660_ (.A1(_0613_),
    .A2(_0621_),
    .B1(_0622_),
    .Y(_0623_));
 sky130_fd_sc_hd__or3_1 _2661_ (.A(_0613_),
    .B(_0622_),
    .C(_0621_),
    .X(_0624_));
 sky130_fd_sc_hd__a31o_1 _2662_ (.A1(_0510_),
    .A2(_0623_),
    .A3(_0624_),
    .B1(_0514_),
    .X(_0625_));
 sky130_fd_sc_hd__o221a_1 _2663_ (.A1(\simon0.play1.tick_counter[12] ),
    .A2(_0570_),
    .B1(_0620_),
    .B2(_0625_),
    .C1(_0618_),
    .X(_0059_));
 sky130_fd_sc_hd__or2b_1 _2664_ (.A(_0619_),
    .B_N(_0443_),
    .X(_0626_));
 sky130_fd_sc_hd__xor2_1 _2665_ (.A(_0445_),
    .B(_0273_),
    .X(_0627_));
 sky130_fd_sc_hd__nand3_1 _2666_ (.A(\simon0.play1.tick_counter[13] ),
    .B(\simon0.play1.tick_counter[12] ),
    .C(_0606_),
    .Y(_0628_));
 sky130_fd_sc_hd__a21o_1 _2667_ (.A1(\simon0.play1.tick_counter[12] ),
    .A2(_0606_),
    .B1(\simon0.play1.tick_counter[13] ),
    .X(_0629_));
 sky130_fd_sc_hd__nand2_1 _2668_ (.A(_0628_),
    .B(_0629_),
    .Y(_0630_));
 sky130_fd_sc_hd__inv_2 _2669_ (.A(_0630_),
    .Y(_0631_));
 sky130_fd_sc_hd__nand2_1 _2670_ (.A(_0627_),
    .B(_0631_),
    .Y(_0632_));
 sky130_fd_sc_hd__nand2_1 _2671_ (.A(_0446_),
    .B(_0630_),
    .Y(_0633_));
 sky130_fd_sc_hd__and2_1 _2672_ (.A(_0632_),
    .B(_0633_),
    .X(_0634_));
 sky130_fd_sc_hd__and3_1 _2673_ (.A(_0626_),
    .B(_0623_),
    .C(_0634_),
    .X(_0635_));
 sky130_fd_sc_hd__a21oi_1 _2674_ (.A1(_0626_),
    .A2(_0623_),
    .B1(_0634_),
    .Y(_0636_));
 sky130_fd_sc_hd__o21a_1 _2675_ (.A1(_0635_),
    .A2(_0636_),
    .B1(_0510_),
    .X(_0637_));
 sky130_fd_sc_hd__a21o_1 _2676_ (.A1(_0489_),
    .A2(_0631_),
    .B1(_0529_),
    .X(_0638_));
 sky130_fd_sc_hd__o221a_1 _2677_ (.A1(\simon0.play1.tick_counter[13] ),
    .A2(_0570_),
    .B1(_0637_),
    .B2(_0638_),
    .C1(_0618_),
    .X(_0060_));
 sky130_fd_sc_hd__nor2_1 _2678_ (.A(_0440_),
    .B(_0628_),
    .Y(_0639_));
 sky130_fd_sc_hd__and2_1 _2679_ (.A(_0440_),
    .B(_0628_),
    .X(_0640_));
 sky130_fd_sc_hd__or2_1 _2680_ (.A(_0639_),
    .B(_0640_),
    .X(_0641_));
 sky130_fd_sc_hd__or2_1 _2681_ (.A(_0501_),
    .B(_0641_),
    .X(_0642_));
 sky130_fd_sc_hd__inv_2 _2682_ (.A(_0626_),
    .Y(_0643_));
 sky130_fd_sc_hd__inv_2 _2683_ (.A(_0608_),
    .Y(_0644_));
 sky130_fd_sc_hd__a221o_1 _2684_ (.A1(_0599_),
    .A2(_0600_),
    .B1(_0644_),
    .B2(_0421_),
    .C1(_0610_),
    .X(_0645_));
 sky130_fd_sc_hd__a32o_1 _2685_ (.A1(_0614_),
    .A2(_0622_),
    .A3(_0645_),
    .B1(_0631_),
    .B2(_0627_),
    .X(_0646_));
 sky130_fd_sc_hd__xor2_1 _2686_ (.A(_0439_),
    .B(_0641_),
    .X(_0647_));
 sky130_fd_sc_hd__o211a_1 _2687_ (.A1(_0643_),
    .A2(_0646_),
    .B1(_0647_),
    .C1(_0633_),
    .X(_0648_));
 sky130_fd_sc_hd__or2_1 _2688_ (.A(_0643_),
    .B(_0646_),
    .X(_0649_));
 sky130_fd_sc_hd__a21oi_1 _2689_ (.A1(_0633_),
    .A2(_0649_),
    .B1(_0647_),
    .Y(_0650_));
 sky130_fd_sc_hd__o31a_1 _2690_ (.A1(_0488_),
    .A2(_0648_),
    .A3(_0650_),
    .B1(_1301_),
    .X(_0651_));
 sky130_fd_sc_hd__a221oi_1 _2691_ (.A1(_0440_),
    .A2(_0529_),
    .B1(_0642_),
    .B2(_0651_),
    .C1(_1201_),
    .Y(_0061_));
 sky130_fd_sc_hd__xnor2_1 _2692_ (.A(\simon0.play1.tick_counter[15] ),
    .B(_0639_),
    .Y(_0652_));
 sky130_fd_sc_hd__nor2_1 _2693_ (.A(_0502_),
    .B(_0652_),
    .Y(_0653_));
 sky130_fd_sc_hd__and2_1 _2694_ (.A(_0436_),
    .B(_0437_),
    .X(_0654_));
 sky130_fd_sc_hd__or2_1 _2695_ (.A(_0654_),
    .B(_0652_),
    .X(_0655_));
 sky130_fd_sc_hd__nand2_1 _2696_ (.A(_0654_),
    .B(_0652_),
    .Y(_0656_));
 sky130_fd_sc_hd__nand2_1 _2697_ (.A(_0655_),
    .B(_0656_),
    .Y(_0657_));
 sky130_fd_sc_hd__nor2_1 _2698_ (.A(_0439_),
    .B(_0641_),
    .Y(_0658_));
 sky130_fd_sc_hd__nor2_1 _2699_ (.A(_0658_),
    .B(_0648_),
    .Y(_0659_));
 sky130_fd_sc_hd__xor2_1 _2700_ (.A(_0657_),
    .B(_0659_),
    .X(_0660_));
 sky130_fd_sc_hd__a21o_1 _2701_ (.A1(_0510_),
    .A2(_0660_),
    .B1(_0529_),
    .X(_0661_));
 sky130_fd_sc_hd__o221a_1 _2702_ (.A1(\simon0.play1.tick_counter[15] ),
    .A2(_0570_),
    .B1(_0653_),
    .B2(_0661_),
    .C1(_0618_),
    .X(_0062_));
 sky130_fd_sc_hd__nor2_1 _2703_ (.A(_0654_),
    .B(_0652_),
    .Y(_0662_));
 sky130_fd_sc_hd__and3_1 _2704_ (.A(\simon0.play1.tick_counter[16] ),
    .B(\simon0.play1.tick_counter[15] ),
    .C(_0639_),
    .X(_0663_));
 sky130_fd_sc_hd__a21oi_1 _2705_ (.A1(\simon0.play1.tick_counter[15] ),
    .A2(_0639_),
    .B1(\simon0.play1.tick_counter[16] ),
    .Y(_0664_));
 sky130_fd_sc_hd__or2_1 _2706_ (.A(_0663_),
    .B(_0664_),
    .X(_0665_));
 sky130_fd_sc_hd__xnor2_1 _2707_ (.A(_0462_),
    .B(_0665_),
    .Y(_0666_));
 sky130_fd_sc_hd__o311a_1 _2708_ (.A1(_0658_),
    .A2(_0648_),
    .A3(_0662_),
    .B1(_0656_),
    .C1(_0666_),
    .X(_0667_));
 sky130_fd_sc_hd__nand2_1 _2709_ (.A(_0655_),
    .B(_0659_),
    .Y(_0668_));
 sky130_fd_sc_hd__a21oi_1 _2710_ (.A1(_0656_),
    .A2(_0668_),
    .B1(_0666_),
    .Y(_0669_));
 sky130_fd_sc_hd__or2_1 _2711_ (.A(_0500_),
    .B(_0665_),
    .X(_0670_));
 sky130_fd_sc_hd__o31a_1 _2712_ (.A1(_0488_),
    .A2(_0667_),
    .A3(_0669_),
    .B1(_0670_),
    .X(_0671_));
 sky130_fd_sc_hd__nand2_1 _2713_ (.A(_0595_),
    .B(_0671_),
    .Y(_0672_));
 sky130_fd_sc_hd__o211a_1 _2714_ (.A1(\simon0.play1.tick_counter[16] ),
    .A2(_1303_),
    .B1(_0672_),
    .C1(_1190_),
    .X(_0063_));
 sky130_fd_sc_hd__xnor2_1 _2715_ (.A(\simon0.play1.tick_counter[17] ),
    .B(_0663_),
    .Y(_0673_));
 sky130_fd_sc_hd__nor2_1 _2716_ (.A(_0502_),
    .B(_0673_),
    .Y(_0674_));
 sky130_fd_sc_hd__nand2_1 _2717_ (.A(_0465_),
    .B(_0466_),
    .Y(_0675_));
 sky130_fd_sc_hd__nor2_1 _2718_ (.A(_0675_),
    .B(_0673_),
    .Y(_0676_));
 sky130_fd_sc_hd__nand2_1 _2719_ (.A(_0675_),
    .B(_0673_),
    .Y(_0677_));
 sky130_fd_sc_hd__or2b_1 _2720_ (.A(_0676_),
    .B_N(_0677_),
    .X(_0678_));
 sky130_fd_sc_hd__or2b_1 _2721_ (.A(_0665_),
    .B_N(_0462_),
    .X(_0679_));
 sky130_fd_sc_hd__inv_2 _2722_ (.A(_0679_),
    .Y(_0680_));
 sky130_fd_sc_hd__or2_1 _2723_ (.A(_0680_),
    .B(_0667_),
    .X(_0681_));
 sky130_fd_sc_hd__xnor2_1 _2724_ (.A(_0678_),
    .B(_0681_),
    .Y(_0682_));
 sky130_fd_sc_hd__a21o_1 _2725_ (.A1(_0510_),
    .A2(_0682_),
    .B1(_0514_),
    .X(_0683_));
 sky130_fd_sc_hd__o221a_1 _2726_ (.A1(\simon0.play1.tick_counter[17] ),
    .A2(_0570_),
    .B1(_0674_),
    .B2(_0683_),
    .C1(_0618_),
    .X(_0064_));
 sky130_fd_sc_hd__and4_1 _2727_ (.A(\simon0.play1.tick_counter[17] ),
    .B(\simon0.play1.tick_counter[16] ),
    .C(\simon0.play1.tick_counter[15] ),
    .D(_0639_),
    .X(_0684_));
 sky130_fd_sc_hd__nor2_1 _2728_ (.A(\simon0.play1.tick_counter[18] ),
    .B(_0684_),
    .Y(_0685_));
 sky130_fd_sc_hd__and2_1 _2729_ (.A(\simon0.play1.tick_counter[18] ),
    .B(_0684_),
    .X(_0686_));
 sky130_fd_sc_hd__or2_1 _2730_ (.A(_0685_),
    .B(_0686_),
    .X(_0687_));
 sky130_fd_sc_hd__xor2_1 _2731_ (.A(_0467_),
    .B(_0687_),
    .X(_0688_));
 sky130_fd_sc_hd__inv_2 _2732_ (.A(_0688_),
    .Y(_0689_));
 sky130_fd_sc_hd__o311a_1 _2733_ (.A1(_0680_),
    .A2(_0667_),
    .A3(_0676_),
    .B1(_0677_),
    .C1(_0689_),
    .X(_0690_));
 sky130_fd_sc_hd__o21a_1 _2734_ (.A1(_0676_),
    .A2(_0681_),
    .B1(_0677_),
    .X(_0691_));
 sky130_fd_sc_hd__nor2_1 _2735_ (.A(_0689_),
    .B(_0691_),
    .Y(_0692_));
 sky130_fd_sc_hd__o31a_1 _2736_ (.A1(_0488_),
    .A2(_0690_),
    .A3(_0692_),
    .B1(_1301_),
    .X(_0693_));
 sky130_fd_sc_hd__o21ai_1 _2737_ (.A1(_0502_),
    .A2(_0687_),
    .B1(_0693_),
    .Y(_0694_));
 sky130_fd_sc_hd__o211a_1 _2738_ (.A1(\simon0.play1.tick_counter[18] ),
    .A2(_1303_),
    .B1(_0694_),
    .C1(_1190_),
    .X(_0065_));
 sky130_fd_sc_hd__xnor2_1 _2739_ (.A(\simon0.play1.tick_counter[19] ),
    .B(_0686_),
    .Y(_0695_));
 sky130_fd_sc_hd__nor2_1 _2740_ (.A(_0510_),
    .B(_0695_),
    .Y(_0696_));
 sky130_fd_sc_hd__and2b_1 _2741_ (.A_N(_0687_),
    .B(_0467_),
    .X(_0697_));
 sky130_fd_sc_hd__or2_1 _2742_ (.A(_0697_),
    .B(_0690_),
    .X(_0698_));
 sky130_fd_sc_hd__nor2_1 _2743_ (.A(_0460_),
    .B(_0695_),
    .Y(_0699_));
 sky130_fd_sc_hd__nand2_1 _2744_ (.A(_0460_),
    .B(_0695_),
    .Y(_0700_));
 sky130_fd_sc_hd__and2b_1 _2745_ (.A_N(_0699_),
    .B(_0700_),
    .X(_0701_));
 sky130_fd_sc_hd__nand2_1 _2746_ (.A(_0698_),
    .B(_0701_),
    .Y(_0702_));
 sky130_fd_sc_hd__or2_1 _2747_ (.A(_0698_),
    .B(_0701_),
    .X(_0703_));
 sky130_fd_sc_hd__a31o_1 _2748_ (.A1(_0510_),
    .A2(_0702_),
    .A3(_0703_),
    .B1(_0514_),
    .X(_0704_));
 sky130_fd_sc_hd__o221a_1 _2749_ (.A1(\simon0.play1.tick_counter[19] ),
    .A2(_0570_),
    .B1(_0696_),
    .B2(_0704_),
    .C1(_0618_),
    .X(_0066_));
 sky130_fd_sc_hd__a21oi_1 _2750_ (.A1(\simon0.play1.tick_counter[19] ),
    .A2(_0686_),
    .B1(\simon0.play1.tick_counter[20] ),
    .Y(_0705_));
 sky130_fd_sc_hd__and3_1 _2751_ (.A(\simon0.play1.tick_counter[20] ),
    .B(\simon0.play1.tick_counter[19] ),
    .C(_0686_),
    .X(_0706_));
 sky130_fd_sc_hd__or2_1 _2752_ (.A(_0705_),
    .B(_0706_),
    .X(_0707_));
 sky130_fd_sc_hd__inv_2 _2753_ (.A(_0707_),
    .Y(_0708_));
 sky130_fd_sc_hd__and2_1 _2754_ (.A(_0392_),
    .B(_0708_),
    .X(_0709_));
 sky130_fd_sc_hd__nor2_1 _2755_ (.A(_0392_),
    .B(_0708_),
    .Y(_0710_));
 sky130_fd_sc_hd__nor2_1 _2756_ (.A(_0709_),
    .B(_0710_),
    .Y(_0711_));
 sky130_fd_sc_hd__a21o_1 _2757_ (.A1(_0698_),
    .A2(_0700_),
    .B1(_0699_),
    .X(_0712_));
 sky130_fd_sc_hd__xnor2_1 _2758_ (.A(_0711_),
    .B(_0712_),
    .Y(_0713_));
 sky130_fd_sc_hd__nor2_1 _2759_ (.A(_0489_),
    .B(_0713_),
    .Y(_0714_));
 sky130_fd_sc_hd__a21o_1 _2760_ (.A1(_0489_),
    .A2(_0708_),
    .B1(_0514_),
    .X(_0715_));
 sky130_fd_sc_hd__o221a_1 _2761_ (.A1(\simon0.play1.tick_counter[20] ),
    .A2(_0570_),
    .B1(_0714_),
    .B2(_0715_),
    .C1(_0618_),
    .X(_0067_));
 sky130_fd_sc_hd__xnor2_2 _2762_ (.A(\simon0.play1.tick_counter[21] ),
    .B(_0706_),
    .Y(_0716_));
 sky130_fd_sc_hd__xor2_1 _2763_ (.A(_0395_),
    .B(_0716_),
    .X(_0717_));
 sky130_fd_sc_hd__a21o_1 _2764_ (.A1(_0711_),
    .A2(_0712_),
    .B1(_0709_),
    .X(_0718_));
 sky130_fd_sc_hd__xnor2_1 _2765_ (.A(_0717_),
    .B(_0718_),
    .Y(_0719_));
 sky130_fd_sc_hd__mux2_1 _2766_ (.A0(_0716_),
    .A1(_0719_),
    .S(_0501_),
    .X(_0720_));
 sky130_fd_sc_hd__nand2_1 _2767_ (.A(_0595_),
    .B(_0720_),
    .Y(_0721_));
 sky130_fd_sc_hd__o211a_1 _2768_ (.A1(\simon0.play1.tick_counter[21] ),
    .A2(_1303_),
    .B1(_0721_),
    .C1(_1190_),
    .X(_0068_));
 sky130_fd_sc_hd__a21oi_1 _2769_ (.A1(\simon0.play1.tick_counter[21] ),
    .A2(_0706_),
    .B1(\simon0.play1.tick_counter[22] ),
    .Y(_0722_));
 sky130_fd_sc_hd__and3_1 _2770_ (.A(\simon0.play1.tick_counter[22] ),
    .B(\simon0.play1.tick_counter[21] ),
    .C(_0706_),
    .X(_0723_));
 sky130_fd_sc_hd__or2_1 _2771_ (.A(_0722_),
    .B(_0723_),
    .X(_0724_));
 sky130_fd_sc_hd__nor2_1 _2772_ (.A(_0389_),
    .B(_0724_),
    .Y(_0725_));
 sky130_fd_sc_hd__nand2_1 _2773_ (.A(_0389_),
    .B(_0724_),
    .Y(_0726_));
 sky130_fd_sc_hd__or2b_1 _2774_ (.A(_0725_),
    .B_N(_0726_),
    .X(_0727_));
 sky130_fd_sc_hd__nor2_1 _2775_ (.A(_0395_),
    .B(_0716_),
    .Y(_0728_));
 sky130_fd_sc_hd__and4_1 _2776_ (.A(_0690_),
    .B(_0701_),
    .C(_0711_),
    .D(_0717_),
    .X(_0729_));
 sky130_fd_sc_hd__a21o_1 _2777_ (.A1(_0697_),
    .A2(_0700_),
    .B1(_0699_),
    .X(_0730_));
 sky130_fd_sc_hd__nand2_1 _2778_ (.A(_0395_),
    .B(_0716_),
    .Y(_0731_));
 sky130_fd_sc_hd__a32o_1 _2779_ (.A1(_0711_),
    .A2(_0717_),
    .A3(_0730_),
    .B1(_0731_),
    .B2(_0709_),
    .X(_0732_));
 sky130_fd_sc_hd__or3_1 _2780_ (.A(_0728_),
    .B(_0729_),
    .C(_0732_),
    .X(_0733_));
 sky130_fd_sc_hd__xor2_1 _2781_ (.A(_0727_),
    .B(_0733_),
    .X(_0734_));
 sky130_fd_sc_hd__mux2_1 _2782_ (.A0(_0724_),
    .A1(_0734_),
    .S(_0501_),
    .X(_0735_));
 sky130_fd_sc_hd__nand2_1 _2783_ (.A(_0595_),
    .B(_0735_),
    .Y(_0736_));
 sky130_fd_sc_hd__o211a_1 _2784_ (.A1(\simon0.play1.tick_counter[22] ),
    .A2(_1303_),
    .B1(_0736_),
    .C1(_1190_),
    .X(_0069_));
 sky130_fd_sc_hd__xnor2_1 _2785_ (.A(\simon0.play1.tick_counter[23] ),
    .B(_0723_),
    .Y(_0737_));
 sky130_fd_sc_hd__nor2_1 _2786_ (.A(_0510_),
    .B(_0737_),
    .Y(_0738_));
 sky130_fd_sc_hd__or2_1 _2787_ (.A(_0388_),
    .B(_0737_),
    .X(_0739_));
 sky130_fd_sc_hd__nand2_1 _2788_ (.A(_0388_),
    .B(_0737_),
    .Y(_0740_));
 sky130_fd_sc_hd__nand2_1 _2789_ (.A(_0739_),
    .B(_0740_),
    .Y(_0741_));
 sky130_fd_sc_hd__a21oi_2 _2790_ (.A1(_0726_),
    .A2(_0733_),
    .B1(_0725_),
    .Y(_0742_));
 sky130_fd_sc_hd__xnor2_1 _2791_ (.A(_0741_),
    .B(_0742_),
    .Y(_0743_));
 sky130_fd_sc_hd__o21ai_1 _2792_ (.A1(_0489_),
    .A2(_0743_),
    .B1(_1302_),
    .Y(_0744_));
 sky130_fd_sc_hd__o221a_1 _2793_ (.A1(\simon0.play1.tick_counter[23] ),
    .A2(_0570_),
    .B1(_0738_),
    .B2(_0744_),
    .C1(_0618_),
    .X(_0070_));
 sky130_fd_sc_hd__a21oi_1 _2794_ (.A1(\simon0.play1.tick_counter[23] ),
    .A2(_0723_),
    .B1(\simon0.play1.tick_counter[24] ),
    .Y(_0745_));
 sky130_fd_sc_hd__and3_1 _2795_ (.A(\simon0.play1.tick_counter[24] ),
    .B(\simon0.play1.tick_counter[23] ),
    .C(_0723_),
    .X(_0746_));
 sky130_fd_sc_hd__or2_1 _2796_ (.A(_0745_),
    .B(_0746_),
    .X(_0747_));
 sky130_fd_sc_hd__inv_2 _2797_ (.A(_0747_),
    .Y(_0748_));
 sky130_fd_sc_hd__nand2_1 _2798_ (.A(_0385_),
    .B(_0748_),
    .Y(_0749_));
 sky130_fd_sc_hd__or2_1 _2799_ (.A(_0385_),
    .B(_0748_),
    .X(_0750_));
 sky130_fd_sc_hd__nand2_1 _2800_ (.A(_0749_),
    .B(_0750_),
    .Y(_0751_));
 sky130_fd_sc_hd__and2_1 _2801_ (.A(_0388_),
    .B(_0737_),
    .X(_0752_));
 sky130_fd_sc_hd__a21o_1 _2802_ (.A1(_0739_),
    .A2(_0742_),
    .B1(_0752_),
    .X(_0753_));
 sky130_fd_sc_hd__nand2_1 _2803_ (.A(_0751_),
    .B(_0753_),
    .Y(_0754_));
 sky130_fd_sc_hd__a211o_1 _2804_ (.A1(_0739_),
    .A2(_0742_),
    .B1(_0751_),
    .C1(_0752_),
    .X(_0755_));
 sky130_fd_sc_hd__and3_1 _2805_ (.A(_0501_),
    .B(_0754_),
    .C(_0755_),
    .X(_0756_));
 sky130_fd_sc_hd__a21o_1 _2806_ (.A1(_0488_),
    .A2(_0748_),
    .B1(_0514_),
    .X(_0757_));
 sky130_fd_sc_hd__o221a_1 _2807_ (.A1(\simon0.play1.tick_counter[24] ),
    .A2(_0570_),
    .B1(_0756_),
    .B2(_0757_),
    .C1(_0618_),
    .X(_0071_));
 sky130_fd_sc_hd__nor2_1 _2808_ (.A(\simon0.play1.tick_counter[25] ),
    .B(_0746_),
    .Y(_0758_));
 sky130_fd_sc_hd__and2_1 _2809_ (.A(\simon0.play1.tick_counter[25] ),
    .B(_0746_),
    .X(_0759_));
 sky130_fd_sc_hd__or2_1 _2810_ (.A(_0758_),
    .B(_0759_),
    .X(_0760_));
 sky130_fd_sc_hd__and4_1 _2811_ (.A(_0500_),
    .B(_0749_),
    .C(_0755_),
    .D(_0760_),
    .X(_0761_));
 sky130_fd_sc_hd__buf_2 _2812_ (.A(_0761_),
    .X(_0762_));
 sky130_fd_sc_hd__and3_1 _2813_ (.A(_0501_),
    .B(_0749_),
    .C(_0755_),
    .X(_0763_));
 sky130_fd_sc_hd__o21ai_1 _2814_ (.A1(_0760_),
    .A2(_0763_),
    .B1(_1302_),
    .Y(_0764_));
 sky130_fd_sc_hd__o221a_1 _2815_ (.A1(\simon0.play1.tick_counter[25] ),
    .A2(_0595_),
    .B1(_0762_),
    .B2(_0764_),
    .C1(_0618_),
    .X(_0072_));
 sky130_fd_sc_hd__xnor2_1 _2816_ (.A(\simon0.play1.tick_counter[26] ),
    .B(_0759_),
    .Y(_0765_));
 sky130_fd_sc_hd__and2_1 _2817_ (.A(_0762_),
    .B(_0765_),
    .X(_0766_));
 sky130_fd_sc_hd__o21ai_1 _2818_ (.A1(_0762_),
    .A2(_0765_),
    .B1(_1302_),
    .Y(_0767_));
 sky130_fd_sc_hd__o221a_1 _2819_ (.A1(\simon0.play1.tick_counter[26] ),
    .A2(_0595_),
    .B1(_0766_),
    .B2(_0767_),
    .C1(_1194_),
    .X(_0073_));
 sky130_fd_sc_hd__a21oi_1 _2820_ (.A1(\simon0.play1.tick_counter[26] ),
    .A2(_0759_),
    .B1(\simon0.play1.tick_counter[27] ),
    .Y(_0768_));
 sky130_fd_sc_hd__and3_1 _2821_ (.A(\simon0.play1.tick_counter[27] ),
    .B(\simon0.play1.tick_counter[26] ),
    .C(_0759_),
    .X(_0769_));
 sky130_fd_sc_hd__or2_1 _2822_ (.A(_0768_),
    .B(_0769_),
    .X(_0770_));
 sky130_fd_sc_hd__nor2_1 _2823_ (.A(_0766_),
    .B(_0770_),
    .Y(_0771_));
 sky130_fd_sc_hd__and2_1 _2824_ (.A(_0765_),
    .B(_0770_),
    .X(_0772_));
 sky130_fd_sc_hd__a21o_1 _2825_ (.A1(_0762_),
    .A2(_0772_),
    .B1(_0514_),
    .X(_0773_));
 sky130_fd_sc_hd__o221a_1 _2826_ (.A1(\simon0.play1.tick_counter[27] ),
    .A2(_0595_),
    .B1(_0771_),
    .B2(_0773_),
    .C1(_1194_),
    .X(_0074_));
 sky130_fd_sc_hd__nor2_1 _2827_ (.A(\simon0.play1.tick_counter[28] ),
    .B(_0769_),
    .Y(_0774_));
 sky130_fd_sc_hd__and2_1 _2828_ (.A(\simon0.play1.tick_counter[28] ),
    .B(_0769_),
    .X(_0775_));
 sky130_fd_sc_hd__or2_1 _2829_ (.A(_0774_),
    .B(_0775_),
    .X(_0776_));
 sky130_fd_sc_hd__a21oi_1 _2830_ (.A1(_0762_),
    .A2(_0772_),
    .B1(_0776_),
    .Y(_0777_));
 sky130_fd_sc_hd__and2_1 _2831_ (.A(_0772_),
    .B(_0776_),
    .X(_0778_));
 sky130_fd_sc_hd__a21o_1 _2832_ (.A1(_0762_),
    .A2(_0778_),
    .B1(_0514_),
    .X(_0779_));
 sky130_fd_sc_hd__o221a_1 _2833_ (.A1(\simon0.play1.tick_counter[28] ),
    .A2(_0595_),
    .B1(_0777_),
    .B2(_0779_),
    .C1(_1194_),
    .X(_0075_));
 sky130_fd_sc_hd__xnor2_1 _2834_ (.A(\simon0.play1.tick_counter[29] ),
    .B(_0775_),
    .Y(_0780_));
 sky130_fd_sc_hd__a21oi_1 _2835_ (.A1(_0762_),
    .A2(_0778_),
    .B1(_0780_),
    .Y(_0781_));
 sky130_fd_sc_hd__and3_1 _2836_ (.A(_0772_),
    .B(_0776_),
    .C(_0780_),
    .X(_0782_));
 sky130_fd_sc_hd__a21o_1 _2837_ (.A1(_0762_),
    .A2(_0782_),
    .B1(_0514_),
    .X(_0783_));
 sky130_fd_sc_hd__o221a_1 _2838_ (.A1(\simon0.play1.tick_counter[29] ),
    .A2(_0595_),
    .B1(_0781_),
    .B2(_0783_),
    .C1(_1194_),
    .X(_0076_));
 sky130_fd_sc_hd__a21oi_1 _2839_ (.A1(\simon0.play1.tick_counter[29] ),
    .A2(_0775_),
    .B1(\simon0.play1.tick_counter[30] ),
    .Y(_0784_));
 sky130_fd_sc_hd__and3_1 _2840_ (.A(\simon0.play1.tick_counter[30] ),
    .B(\simon0.play1.tick_counter[29] ),
    .C(_0775_),
    .X(_0785_));
 sky130_fd_sc_hd__or2_1 _2841_ (.A(_0784_),
    .B(_0785_),
    .X(_0786_));
 sky130_fd_sc_hd__and3_1 _2842_ (.A(_0762_),
    .B(_0782_),
    .C(_0786_),
    .X(_0787_));
 sky130_fd_sc_hd__a21o_1 _2843_ (.A1(_0762_),
    .A2(_0782_),
    .B1(_0786_),
    .X(_0788_));
 sky130_fd_sc_hd__nand2_1 _2844_ (.A(_1302_),
    .B(_0788_),
    .Y(_0789_));
 sky130_fd_sc_hd__o221a_1 _2845_ (.A1(\simon0.play1.tick_counter[30] ),
    .A2(_0595_),
    .B1(_0787_),
    .B2(_0789_),
    .C1(_1194_),
    .X(_0077_));
 sky130_fd_sc_hd__a21o_1 _2846_ (.A1(_0761_),
    .A2(_0782_),
    .B1(_0785_),
    .X(_0790_));
 sky130_fd_sc_hd__nand3b_1 _2847_ (.A_N(_0784_),
    .B(_0782_),
    .C(_0761_),
    .Y(_0791_));
 sky130_fd_sc_hd__a41o_1 _2848_ (.A1(\simon0.play1.tick_counter[31] ),
    .A2(_1301_),
    .A3(_0790_),
    .A4(_0791_),
    .B1(net4),
    .X(_0792_));
 sky130_fd_sc_hd__a31o_1 _2849_ (.A1(_1301_),
    .A2(_0790_),
    .A3(_0791_),
    .B1(\simon0.play1.tick_counter[31] ),
    .X(_0793_));
 sky130_fd_sc_hd__and2b_1 _2850_ (.A_N(_0792_),
    .B(_0793_),
    .X(_0794_));
 sky130_fd_sc_hd__clkbuf_1 _2851_ (.A(_0794_),
    .X(_0078_));
 sky130_fd_sc_hd__a211oi_1 _2852_ (.A1(\simon0.play1.sound ),
    .A2(_0502_),
    .B1(_0529_),
    .C1(_1123_),
    .Y(_0795_));
 sky130_fd_sc_hd__o21a_1 _2853_ (.A1(\simon0.play1.sound ),
    .A2(_0502_),
    .B1(_0795_),
    .X(_0079_));
 sky130_fd_sc_hd__nand2_1 _2854_ (.A(_1216_),
    .B(_1289_),
    .Y(_0796_));
 sky130_fd_sc_hd__mux2_1 _2855_ (.A0(_1213_),
    .A1(\simon0.seq[20][0] ),
    .S(_0796_),
    .X(_0797_));
 sky130_fd_sc_hd__clkbuf_1 _2856_ (.A(_0797_),
    .X(_0080_));
 sky130_fd_sc_hd__mux2_1 _2857_ (.A0(_1223_),
    .A1(\simon0.seq[20][1] ),
    .S(_0796_),
    .X(_0798_));
 sky130_fd_sc_hd__clkbuf_1 _2858_ (.A(_0798_),
    .X(_0081_));
 sky130_fd_sc_hd__nor2_1 _2859_ (.A(_1124_),
    .B(\simon0.next_random[0] ),
    .Y(_0082_));
 sky130_fd_sc_hd__a21oi_1 _2860_ (.A1(\simon0.next_random[0] ),
    .A2(\simon0.next_random[1] ),
    .B1(_1123_),
    .Y(_0799_));
 sky130_fd_sc_hd__o21a_1 _2861_ (.A1(\simon0.next_random[0] ),
    .A2(\simon0.next_random[1] ),
    .B1(_0799_),
    .X(_0083_));
 sky130_fd_sc_hd__buf_2 _2862_ (.A(\simon0.tone_sequence_counter[2] ),
    .X(_0800_));
 sky130_fd_sc_hd__nor2_2 _2863_ (.A(\simon0.tone_sequence_counter[0] ),
    .B(\simon0.tone_sequence_counter[1] ),
    .Y(_0801_));
 sky130_fd_sc_hd__nand2_2 _2864_ (.A(_0800_),
    .B(_0801_),
    .Y(_0802_));
 sky130_fd_sc_hd__nand2_1 _2865_ (.A(\simon0.millis_counter[8] ),
    .B(\simon0.millis_counter[9] ),
    .Y(_0803_));
 sky130_fd_sc_hd__and3_1 _2866_ (.A(\simon0.millis_counter[3] ),
    .B(\simon0.millis_counter[6] ),
    .C(\simon0.millis_counter[7] ),
    .X(_0804_));
 sky130_fd_sc_hd__or4b_2 _2867_ (.A(_1107_),
    .B(_1172_),
    .C(_0803_),
    .D_N(_0804_),
    .X(_0805_));
 sky130_fd_sc_hd__or2_1 _2868_ (.A(\simon0.tone_sequence_counter[2] ),
    .B(_1173_),
    .X(_0806_));
 sky130_fd_sc_hd__o211a_1 _2869_ (.A1(_0802_),
    .A2(_0805_),
    .B1(\simon0.state[7] ),
    .C1(_0806_),
    .X(_0807_));
 sky130_fd_sc_hd__nor2_2 _2870_ (.A(_1197_),
    .B(_1115_),
    .Y(_0808_));
 sky130_fd_sc_hd__or3_1 _2871_ (.A(\simon0.state[4] ),
    .B(_1112_),
    .C(\simon0.state[7] ),
    .X(_0809_));
 sky130_fd_sc_hd__or4b_2 _2872_ (.A(net4),
    .B(_0807_),
    .C(_0808_),
    .D_N(_0809_),
    .X(_0810_));
 sky130_fd_sc_hd__o21ba_1 _2873_ (.A1(_1112_),
    .A2(\simon0.state[7] ),
    .B1_N(_0810_),
    .X(_0811_));
 sky130_fd_sc_hd__mux2_1 _2874_ (.A0(_0811_),
    .A1(_0810_),
    .S(\simon0.tone_sequence_counter[0] ),
    .X(_0812_));
 sky130_fd_sc_hd__clkbuf_1 _2875_ (.A(_0812_),
    .X(_0084_));
 sky130_fd_sc_hd__and2_1 _2876_ (.A(\simon0.tone_sequence_counter[0] ),
    .B(\simon0.tone_sequence_counter[1] ),
    .X(_0813_));
 sky130_fd_sc_hd__and2_1 _2877_ (.A(_0800_),
    .B(_0801_),
    .X(_0814_));
 sky130_fd_sc_hd__a2bb2o_1 _2878_ (.A1_N(_0813_),
    .A2_N(_0801_),
    .B1(_0814_),
    .B2(\simon0.state[7] ),
    .X(_0815_));
 sky130_fd_sc_hd__a22o_1 _2879_ (.A1(\simon0.tone_sequence_counter[1] ),
    .A2(_0810_),
    .B1(_0811_),
    .B2(_0815_),
    .X(_0085_));
 sky130_fd_sc_hd__nand2_1 _2880_ (.A(_0800_),
    .B(_0813_),
    .Y(_0816_));
 sky130_fd_sc_hd__or2_1 _2881_ (.A(_0800_),
    .B(_0813_),
    .X(_0817_));
 sky130_fd_sc_hd__a32o_1 _2882_ (.A1(_0816_),
    .A2(_0811_),
    .A3(_0817_),
    .B1(_0810_),
    .B2(_0800_),
    .X(_0086_));
 sky130_fd_sc_hd__and3_1 _2883_ (.A(_1187_),
    .B(_0806_),
    .C(_0802_),
    .X(_0818_));
 sky130_fd_sc_hd__and2_1 _2884_ (.A(_1085_),
    .B(_1173_),
    .X(_0819_));
 sky130_fd_sc_hd__nor2_1 _2885_ (.A(\simon0.state[2] ),
    .B(_1205_),
    .Y(_0820_));
 sky130_fd_sc_hd__nor4_4 _2886_ (.A(_0808_),
    .B(_0818_),
    .C(_0819_),
    .D(_0820_),
    .Y(_0821_));
 sky130_fd_sc_hd__buf_2 _2887_ (.A(_0821_),
    .X(_0822_));
 sky130_fd_sc_hd__nor2_1 _2888_ (.A(\simon0.tone_sequence_counter[1] ),
    .B(_0800_),
    .Y(_0823_));
 sky130_fd_sc_hd__and2b_1 _2889_ (.A_N(\simon0.tone_sequence_counter[1] ),
    .B(\simon0.tone_sequence_counter[0] ),
    .X(_0824_));
 sky130_fd_sc_hd__nand2_1 _2890_ (.A(\simon0.tone_sequence_counter[1] ),
    .B(_0800_),
    .Y(_0825_));
 sky130_fd_sc_hd__or3b_1 _2891_ (.A(_0824_),
    .B(_1197_),
    .C_N(_0825_),
    .X(_0826_));
 sky130_fd_sc_hd__nor2_1 _2892_ (.A(\simon0.millis_counter[0] ),
    .B(_0802_),
    .Y(_0827_));
 sky130_fd_sc_hd__a21oi_1 _2893_ (.A1(_0805_),
    .A2(_0827_),
    .B1(\simon0.tone_sequence_counter[0] ),
    .Y(_0828_));
 sky130_fd_sc_hd__nand2_1 _2894_ (.A(\simon0.state[7] ),
    .B(_1184_),
    .Y(_0829_));
 sky130_fd_sc_hd__o221ai_1 _2895_ (.A1(_0823_),
    .A2(_0826_),
    .B1(_0828_),
    .B2(_0829_),
    .C1(_0821_),
    .Y(_0830_));
 sky130_fd_sc_hd__o211a_1 _2896_ (.A1(\simon0.play1.freq[0] ),
    .A2(_0822_),
    .B1(_0830_),
    .C1(_1190_),
    .X(_0087_));
 sky130_fd_sc_hd__or2_1 _2897_ (.A(_1147_),
    .B(_1166_),
    .X(_0831_));
 sky130_fd_sc_hd__nand2_1 _2898_ (.A(_1147_),
    .B(_1166_),
    .Y(_0832_));
 sky130_fd_sc_hd__nand2_1 _2899_ (.A(_0831_),
    .B(_0832_),
    .Y(_0833_));
 sky130_fd_sc_hd__nand2_2 _2900_ (.A(_1169_),
    .B(_1173_),
    .Y(_0834_));
 sky130_fd_sc_hd__nand2_1 _2901_ (.A(\simon0.user_input[0] ),
    .B(\simon0.user_input[1] ),
    .Y(_0835_));
 sky130_fd_sc_hd__or2_1 _2902_ (.A(\simon0.user_input[0] ),
    .B(\simon0.user_input[1] ),
    .X(_0836_));
 sky130_fd_sc_hd__nand2_1 _2903_ (.A(_0835_),
    .B(_0836_),
    .Y(_0837_));
 sky130_fd_sc_hd__nand2_1 _2904_ (.A(\simon0.millis_counter[0] ),
    .B(\simon0.millis_counter[1] ),
    .Y(_0838_));
 sky130_fd_sc_hd__o21ai_1 _2905_ (.A1(_0802_),
    .A2(_0805_),
    .B1(_1187_),
    .Y(_0839_));
 sky130_fd_sc_hd__a31o_1 _2906_ (.A1(_1106_),
    .A2(_0814_),
    .A3(_0838_),
    .B1(_0839_),
    .X(_0840_));
 sky130_fd_sc_hd__o211a_1 _2907_ (.A1(_0834_),
    .A2(_0837_),
    .B1(_0840_),
    .C1(_0826_),
    .X(_0841_));
 sky130_fd_sc_hd__o211a_1 _2908_ (.A1(_1205_),
    .A2(_0833_),
    .B1(_0841_),
    .C1(_0821_),
    .X(_0842_));
 sky130_fd_sc_hd__o21ai_1 _2909_ (.A1(\simon0.play1.freq[1] ),
    .A2(_0821_),
    .B1(_1194_),
    .Y(_0843_));
 sky130_fd_sc_hd__nor2_1 _2910_ (.A(_0842_),
    .B(_0843_),
    .Y(_0088_));
 sky130_fd_sc_hd__inv_2 _2911_ (.A(_0821_),
    .Y(_0844_));
 sky130_fd_sc_hd__nand2_1 _2912_ (.A(\simon0.millis_counter[2] ),
    .B(_1106_),
    .Y(_0845_));
 sky130_fd_sc_hd__a21bo_1 _2913_ (.A1(_1107_),
    .A2(_0845_),
    .B1_N(_0800_),
    .X(_0846_));
 sky130_fd_sc_hd__a32o_1 _2914_ (.A1(_1187_),
    .A2(_0801_),
    .A3(_0846_),
    .B1(_1191_),
    .B2(_1149_),
    .X(_0847_));
 sky130_fd_sc_hd__a21oi_1 _2915_ (.A1(_1157_),
    .A2(_1165_),
    .B1(_1205_),
    .Y(_0848_));
 sky130_fd_sc_hd__or2_1 _2916_ (.A(\simon0.play1.freq[2] ),
    .B(_0821_),
    .X(_0849_));
 sky130_fd_sc_hd__o311a_1 _2917_ (.A1(_0844_),
    .A2(_0847_),
    .A3(_0848_),
    .B1(_0849_),
    .C1(_1194_),
    .X(_0089_));
 sky130_fd_sc_hd__a21o_1 _2918_ (.A1(_1138_),
    .A2(_1146_),
    .B1(_1205_),
    .X(_0850_));
 sky130_fd_sc_hd__or2_1 _2919_ (.A(_1166_),
    .B(_0850_),
    .X(_0851_));
 sky130_fd_sc_hd__a21o_1 _2920_ (.A1(\simon0.millis_counter[2] ),
    .A2(_1106_),
    .B1(\simon0.millis_counter[3] ),
    .X(_0852_));
 sky130_fd_sc_hd__nand3_1 _2921_ (.A(\simon0.millis_counter[2] ),
    .B(\simon0.millis_counter[3] ),
    .C(_1106_),
    .Y(_0853_));
 sky130_fd_sc_hd__a31o_1 _2922_ (.A1(_0814_),
    .A2(_0852_),
    .A3(_0853_),
    .B1(_0829_),
    .X(_0854_));
 sky130_fd_sc_hd__mux2_1 _2923_ (.A0(\simon0.tone_sequence_counter[1] ),
    .A1(_0800_),
    .S(\simon0.tone_sequence_counter[0] ),
    .X(_0855_));
 sky130_fd_sc_hd__o32a_1 _2924_ (.A1(\simon0.user_input[0] ),
    .A2(_1149_),
    .A3(_0834_),
    .B1(_0855_),
    .B2(_1197_),
    .X(_0856_));
 sky130_fd_sc_hd__a41o_1 _2925_ (.A1(_0821_),
    .A2(_0851_),
    .A3(_0854_),
    .A4(_0856_),
    .B1(_1123_),
    .X(_0857_));
 sky130_fd_sc_hd__o21ba_1 _2926_ (.A1(\simon0.play1.freq[3] ),
    .A2(_0822_),
    .B1_N(_0857_),
    .X(_0090_));
 sky130_fd_sc_hd__nor2_1 _2927_ (.A(_1205_),
    .B(_0831_),
    .Y(_0858_));
 sky130_fd_sc_hd__nor2_1 _2928_ (.A(_0829_),
    .B(_0802_),
    .Y(_0859_));
 sky130_fd_sc_hd__and3_1 _2929_ (.A(_1112_),
    .B(_0825_),
    .C(_0855_),
    .X(_0860_));
 sky130_fd_sc_hd__a31o_1 _2930_ (.A1(\simon0.millis_counter[4] ),
    .A2(_0852_),
    .A3(_0859_),
    .B1(_0860_),
    .X(_0861_));
 sky130_fd_sc_hd__nor2_1 _2931_ (.A(_0834_),
    .B(_0835_),
    .Y(_0862_));
 sky130_fd_sc_hd__or2_1 _2932_ (.A(\simon0.millis_counter[4] ),
    .B(_0852_),
    .X(_0863_));
 sky130_fd_sc_hd__or3_1 _2933_ (.A(_0829_),
    .B(_0802_),
    .C(_0863_),
    .X(_0864_));
 sky130_fd_sc_hd__or4b_1 _2934_ (.A(_0844_),
    .B(_0861_),
    .C(_0862_),
    .D_N(_0864_),
    .X(_0865_));
 sky130_fd_sc_hd__o221a_1 _2935_ (.A1(\simon0.play1.freq[4] ),
    .A2(_0822_),
    .B1(_0858_),
    .B2(_0865_),
    .C1(_1194_),
    .X(_0091_));
 sky130_fd_sc_hd__a21o_1 _2936_ (.A1(_0814_),
    .A2(_0863_),
    .B1(_0829_),
    .X(_0866_));
 sky130_fd_sc_hd__o21ai_1 _2937_ (.A1(\simon0.tone_sequence_counter[0] ),
    .A2(_0866_),
    .B1(_0822_),
    .Y(_0867_));
 sky130_fd_sc_hd__o211a_1 _2938_ (.A1(\simon0.play1.freq[5] ),
    .A2(_0822_),
    .B1(_0867_),
    .C1(_0499_),
    .X(_0092_));
 sky130_fd_sc_hd__nand2_1 _2939_ (.A(_1112_),
    .B(_0801_),
    .Y(_0868_));
 sky130_fd_sc_hd__o221a_1 _2940_ (.A1(\simon0.user_input[0] ),
    .A2(_0834_),
    .B1(_0866_),
    .B2(\simon0.tone_sequence_counter[1] ),
    .C1(_0868_),
    .X(_0869_));
 sky130_fd_sc_hd__a31o_1 _2941_ (.A1(_0821_),
    .A2(_0850_),
    .A3(_0869_),
    .B1(_1123_),
    .X(_0870_));
 sky130_fd_sc_hd__o21ba_1 _2942_ (.A1(\simon0.play1.freq[6] ),
    .A2(_0822_),
    .B1_N(_0870_),
    .X(_0093_));
 sky130_fd_sc_hd__a21o_1 _2943_ (.A1(_1147_),
    .A2(_1166_),
    .B1(_1205_),
    .X(_0871_));
 sky130_fd_sc_hd__inv_2 _2944_ (.A(_0871_),
    .Y(_0872_));
 sky130_fd_sc_hd__o31a_1 _2945_ (.A1(_1197_),
    .A2(_0801_),
    .A3(_0817_),
    .B1(_1205_),
    .X(_0873_));
 sky130_fd_sc_hd__o311a_1 _2946_ (.A1(\simon0.user_input[0] ),
    .A2(\simon0.user_input[1] ),
    .A3(_0834_),
    .B1(_0864_),
    .C1(_0873_),
    .X(_0874_));
 sky130_fd_sc_hd__o21ai_1 _2947_ (.A1(_0872_),
    .A2(_0874_),
    .B1(_0822_),
    .Y(_0875_));
 sky130_fd_sc_hd__o211a_1 _2948_ (.A1(\simon0.play1.freq[7] ),
    .A2(_0822_),
    .B1(_0875_),
    .C1(_0499_),
    .X(_0094_));
 sky130_fd_sc_hd__or2_1 _2949_ (.A(_0824_),
    .B(_0823_),
    .X(_0876_));
 sky130_fd_sc_hd__a22o_1 _2950_ (.A1(_1112_),
    .A2(_0876_),
    .B1(_0836_),
    .B2(_1191_),
    .X(_0877_));
 sky130_fd_sc_hd__or3b_1 _2951_ (.A(_0844_),
    .B(_0877_),
    .C_N(_0864_),
    .X(_0878_));
 sky130_fd_sc_hd__o221a_1 _2952_ (.A1(\simon0.play1.freq[8] ),
    .A2(_0822_),
    .B1(_0872_),
    .B2(_0878_),
    .C1(_1194_),
    .X(_0095_));
 sky130_fd_sc_hd__o21ba_1 _2953_ (.A1(_0802_),
    .A2(_0863_),
    .B1_N(_0839_),
    .X(_0879_));
 sky130_fd_sc_hd__or2_1 _2954_ (.A(\simon0.tone_sequence_counter[1] ),
    .B(_0800_),
    .X(_0880_));
 sky130_fd_sc_hd__a31o_1 _2955_ (.A1(_1112_),
    .A2(_0825_),
    .A3(_0880_),
    .B1(_0862_),
    .X(_0881_));
 sky130_fd_sc_hd__or4_1 _2956_ (.A(_0844_),
    .B(_0858_),
    .C(_0879_),
    .D(_0881_),
    .X(_0882_));
 sky130_fd_sc_hd__o211a_1 _2957_ (.A1(\simon0.play1.freq[9] ),
    .A2(_0822_),
    .B1(_0882_),
    .C1(_0499_),
    .X(_0096_));
 sky130_fd_sc_hd__xnor2_1 _2958_ (.A(\simon0.tick_counter[14] ),
    .B(_1337_),
    .Y(_0883_));
 sky130_fd_sc_hd__a2bb2o_1 _2959_ (.A1_N(\simon0.tick_counter[7] ),
    .A2_N(_1434_),
    .B1(_1312_),
    .B2(\simon0.tick_counter[13] ),
    .X(_0884_));
 sky130_fd_sc_hd__a2bb2o_1 _2960_ (.A1_N(\simon0.tick_counter[4] ),
    .A2_N(_0191_),
    .B1(_0398_),
    .B2(\simon0.tick_counter[1] ),
    .X(_0885_));
 sky130_fd_sc_hd__xnor2_1 _2961_ (.A(\simon0.tick_counter[6] ),
    .B(_1420_),
    .Y(_0886_));
 sky130_fd_sc_hd__or4_1 _2962_ (.A(_0883_),
    .B(_0884_),
    .C(_0885_),
    .D(_0886_),
    .X(_0887_));
 sky130_fd_sc_hd__o22ai_1 _2963_ (.A1(\simon0.tick_counter[9] ),
    .A2(_1367_),
    .B1(_1395_),
    .B2(\simon0.tick_counter[8] ),
    .Y(_0888_));
 sky130_fd_sc_hd__a22o_1 _2964_ (.A1(\simon0.tick_counter[15] ),
    .A2(_1308_),
    .B1(_1395_),
    .B2(\simon0.tick_counter[8] ),
    .X(_0889_));
 sky130_fd_sc_hd__a2bb2o_1 _2965_ (.A1_N(\simon0.tick_counter[15] ),
    .A2_N(_1308_),
    .B1(_1434_),
    .B2(\simon0.tick_counter[7] ),
    .X(_0890_));
 sky130_fd_sc_hd__a221o_1 _2966_ (.A1(\simon0.tick_counter[0] ),
    .A2(_0242_),
    .B1(_0243_),
    .B2(\simon0.tick_counter[2] ),
    .C1(_0890_),
    .X(_0891_));
 sky130_fd_sc_hd__or4_1 _2967_ (.A(_0887_),
    .B(_0888_),
    .C(_0889_),
    .D(_0891_),
    .X(_0892_));
 sky130_fd_sc_hd__or2_1 _2968_ (.A(\simon0.tick_counter[1] ),
    .B(_0398_),
    .X(_0893_));
 sky130_fd_sc_hd__a22o_1 _2969_ (.A1(\simon0.tick_counter[9] ),
    .A2(_1367_),
    .B1(_0195_),
    .B2(\simon0.tick_counter[3] ),
    .X(_0894_));
 sky130_fd_sc_hd__xnor2_1 _2970_ (.A(\simon0.tick_counter[11] ),
    .B(_1315_),
    .Y(_0895_));
 sky130_fd_sc_hd__o2bb2a_1 _2971_ (.A1_N(\simon0.tick_counter[4] ),
    .A2_N(_0191_),
    .B1(_1320_),
    .B2(\simon0.tick_counter[12] ),
    .X(_0896_));
 sky130_fd_sc_hd__o22a_1 _2972_ (.A1(\simon0.tick_counter[3] ),
    .A2(_0195_),
    .B1(_0243_),
    .B2(\simon0.tick_counter[2] ),
    .X(_0897_));
 sky130_fd_sc_hd__and4b_1 _2973_ (.A_N(_0894_),
    .B(_0895_),
    .C(_0896_),
    .D(_0897_),
    .X(_0898_));
 sky130_fd_sc_hd__xnor2_1 _2974_ (.A(\simon0.tick_counter[5] ),
    .B(_1426_),
    .Y(_0899_));
 sky130_fd_sc_hd__o2bb2a_1 _2975_ (.A1_N(\simon0.tick_counter[12] ),
    .A2_N(_1320_),
    .B1(_0242_),
    .B2(\simon0.tick_counter[0] ),
    .X(_0900_));
 sky130_fd_sc_hd__xnor2_1 _2976_ (.A(\simon0.tick_counter[10] ),
    .B(_1329_),
    .Y(_0901_));
 sky130_fd_sc_hd__o2111a_1 _2977_ (.A1(\simon0.tick_counter[13] ),
    .A2(_1312_),
    .B1(_0899_),
    .C1(_0900_),
    .D1(_0901_),
    .X(_0902_));
 sky130_fd_sc_hd__and4b_1 _2978_ (.A_N(_0892_),
    .B(_0893_),
    .C(_0898_),
    .D(_0902_),
    .X(_0903_));
 sky130_fd_sc_hd__buf_2 _2979_ (.A(_0903_),
    .X(_0904_));
 sky130_fd_sc_hd__a21oi_1 _2980_ (.A1(\simon0.millis_counter[0] ),
    .A2(_0904_),
    .B1(_1123_),
    .Y(_0905_));
 sky130_fd_sc_hd__a21o_1 _2981_ (.A1(\simon0.state[0] ),
    .A2(_1184_),
    .B1(_1206_),
    .X(_0906_));
 sky130_fd_sc_hd__a211o_1 _2982_ (.A1(_1173_),
    .A2(_1187_),
    .B1(_0859_),
    .C1(_0906_),
    .X(_0907_));
 sky130_fd_sc_hd__a211o_1 _2983_ (.A1(_1169_),
    .A2(_1168_),
    .B1(_1191_),
    .C1(_0907_),
    .X(_0908_));
 sky130_fd_sc_hd__o21ai_1 _2984_ (.A1(_1104_),
    .A2(_1110_),
    .B1(_1085_),
    .Y(_0909_));
 sky130_fd_sc_hd__or3b_1 _2985_ (.A(_0808_),
    .B(_0908_),
    .C_N(_0909_),
    .X(_0910_));
 sky130_fd_sc_hd__o211a_1 _2986_ (.A1(\simon0.millis_counter[0] ),
    .A2(_0904_),
    .B1(_0905_),
    .C1(_0910_),
    .X(_0097_));
 sky130_fd_sc_hd__a21oi_1 _2987_ (.A1(\simon0.millis_counter[0] ),
    .A2(_0904_),
    .B1(\simon0.millis_counter[1] ),
    .Y(_0911_));
 sky130_fd_sc_hd__or4_1 _2988_ (.A(_1169_),
    .B(_1187_),
    .C(_0808_),
    .D(_0906_),
    .X(_0912_));
 sky130_fd_sc_hd__nor2_1 _2989_ (.A(_1085_),
    .B(_0912_),
    .Y(_0913_));
 sky130_fd_sc_hd__and3_1 _2990_ (.A(\simon0.millis_counter[0] ),
    .B(\simon0.millis_counter[1] ),
    .C(_0904_),
    .X(_0914_));
 sky130_fd_sc_hd__nor4_1 _2991_ (.A(_1123_),
    .B(_0911_),
    .C(_0913_),
    .D(_0914_),
    .Y(_0098_));
 sky130_fd_sc_hd__nor3_1 _2992_ (.A(_1085_),
    .B(_0808_),
    .C(_0908_),
    .Y(_0915_));
 sky130_fd_sc_hd__nor2_1 _2993_ (.A(\simon0.millis_counter[2] ),
    .B(_0914_),
    .Y(_0916_));
 sky130_fd_sc_hd__and2_1 _2994_ (.A(\simon0.millis_counter[2] ),
    .B(_0914_),
    .X(_0917_));
 sky130_fd_sc_hd__nor4_1 _2995_ (.A(_1123_),
    .B(_0915_),
    .C(_0916_),
    .D(_0917_),
    .Y(_0099_));
 sky130_fd_sc_hd__o31a_1 _2996_ (.A1(_1085_),
    .A2(_1112_),
    .A3(_0908_),
    .B1(_1084_),
    .X(_0918_));
 sky130_fd_sc_hd__o21ai_1 _2997_ (.A1(\simon0.millis_counter[3] ),
    .A2(_0917_),
    .B1(_0918_),
    .Y(_0919_));
 sky130_fd_sc_hd__and3_1 _2998_ (.A(\simon0.millis_counter[2] ),
    .B(\simon0.millis_counter[3] ),
    .C(_0914_),
    .X(_0920_));
 sky130_fd_sc_hd__nor2_1 _2999_ (.A(_0919_),
    .B(_0920_),
    .Y(_0100_));
 sky130_fd_sc_hd__inv_2 _3000_ (.A(_0912_),
    .Y(_0921_));
 sky130_fd_sc_hd__a21oi_1 _3001_ (.A1(_0909_),
    .A2(_0921_),
    .B1(net4),
    .Y(_0922_));
 sky130_fd_sc_hd__or2_1 _3002_ (.A(\simon0.millis_counter[4] ),
    .B(_0920_),
    .X(_0923_));
 sky130_fd_sc_hd__nand2_1 _3003_ (.A(\simon0.millis_counter[4] ),
    .B(_0920_),
    .Y(_0924_));
 sky130_fd_sc_hd__and3_1 _3004_ (.A(_0922_),
    .B(_0923_),
    .C(_0924_),
    .X(_0925_));
 sky130_fd_sc_hd__clkbuf_1 _3005_ (.A(_0925_),
    .X(_0101_));
 sky130_fd_sc_hd__and3_1 _3006_ (.A(\simon0.millis_counter[4] ),
    .B(\simon0.millis_counter[5] ),
    .C(_0920_),
    .X(_0926_));
 sky130_fd_sc_hd__a21o_1 _3007_ (.A1(\simon0.millis_counter[4] ),
    .A2(_0920_),
    .B1(\simon0.millis_counter[5] ),
    .X(_0927_));
 sky130_fd_sc_hd__and3b_1 _3008_ (.A_N(_0926_),
    .B(_0918_),
    .C(_0927_),
    .X(_0928_));
 sky130_fd_sc_hd__clkbuf_1 _3009_ (.A(_0928_),
    .X(_0102_));
 sky130_fd_sc_hd__or2_1 _3010_ (.A(\simon0.millis_counter[6] ),
    .B(_0926_),
    .X(_0929_));
 sky130_fd_sc_hd__o31a_1 _3011_ (.A1(_1187_),
    .A2(_1203_),
    .A3(_0906_),
    .B1(_1084_),
    .X(_0930_));
 sky130_fd_sc_hd__nand2_1 _3012_ (.A(\simon0.millis_counter[6] ),
    .B(_0926_),
    .Y(_0931_));
 sky130_fd_sc_hd__and3_1 _3013_ (.A(_0929_),
    .B(_0930_),
    .C(_0931_),
    .X(_0932_));
 sky130_fd_sc_hd__clkbuf_1 _3014_ (.A(_0932_),
    .X(_0103_));
 sky130_fd_sc_hd__a21o_1 _3015_ (.A1(\simon0.millis_counter[6] ),
    .A2(_0926_),
    .B1(\simon0.millis_counter[7] ),
    .X(_0933_));
 sky130_fd_sc_hd__nand3_1 _3016_ (.A(\simon0.millis_counter[6] ),
    .B(\simon0.millis_counter[7] ),
    .C(_0926_),
    .Y(_0934_));
 sky130_fd_sc_hd__and3_1 _3017_ (.A(_0922_),
    .B(_0933_),
    .C(_0934_),
    .X(_0935_));
 sky130_fd_sc_hd__clkbuf_1 _3018_ (.A(_0935_),
    .X(_0104_));
 sky130_fd_sc_hd__or4_1 _3019_ (.A(_1112_),
    .B(_1189_),
    .C(_1191_),
    .D(_0907_),
    .X(_0936_));
 sky130_fd_sc_hd__xnor2_1 _3020_ (.A(\simon0.millis_counter[8] ),
    .B(_0934_),
    .Y(_0937_));
 sky130_fd_sc_hd__a21bo_1 _3021_ (.A1(_1085_),
    .A2(_1111_),
    .B1_N(_1199_),
    .X(_0938_));
 sky130_fd_sc_hd__a22o_1 _3022_ (.A1(_0936_),
    .A2(_0937_),
    .B1(_0938_),
    .B2(_1104_),
    .X(_0939_));
 sky130_fd_sc_hd__and2_1 _3023_ (.A(_1084_),
    .B(_0939_),
    .X(_0940_));
 sky130_fd_sc_hd__clkbuf_1 _3024_ (.A(_0940_),
    .X(_0105_));
 sky130_fd_sc_hd__and3_1 _3025_ (.A(\simon0.millis_counter[6] ),
    .B(\simon0.millis_counter[7] ),
    .C(_0926_),
    .X(_0941_));
 sky130_fd_sc_hd__a21o_1 _3026_ (.A1(\simon0.millis_counter[8] ),
    .A2(_0941_),
    .B1(\simon0.millis_counter[9] ),
    .X(_0942_));
 sky130_fd_sc_hd__o211a_1 _3027_ (.A1(_0803_),
    .A2(_0934_),
    .B1(_0942_),
    .C1(_0930_),
    .X(_0106_));
 sky130_fd_sc_hd__nor2_2 _3028_ (.A(net4),
    .B(_0904_),
    .Y(_0943_));
 sky130_fd_sc_hd__buf_2 _3029_ (.A(_0943_),
    .X(_0944_));
 sky130_fd_sc_hd__and2b_1 _3030_ (.A_N(\simon0.tick_counter[0] ),
    .B(_0944_),
    .X(_0945_));
 sky130_fd_sc_hd__clkbuf_1 _3031_ (.A(_0945_),
    .X(_0107_));
 sky130_fd_sc_hd__a21boi_1 _3032_ (.A1(\simon0.tick_counter[1] ),
    .A2(\simon0.tick_counter[0] ),
    .B1_N(_0944_),
    .Y(_0946_));
 sky130_fd_sc_hd__o21a_1 _3033_ (.A1(\simon0.tick_counter[1] ),
    .A2(\simon0.tick_counter[0] ),
    .B1(_0946_),
    .X(_0108_));
 sky130_fd_sc_hd__and3_1 _3034_ (.A(\simon0.tick_counter[1] ),
    .B(\simon0.tick_counter[0] ),
    .C(\simon0.tick_counter[2] ),
    .X(_0947_));
 sky130_fd_sc_hd__a21o_1 _3035_ (.A1(\simon0.tick_counter[1] ),
    .A2(\simon0.tick_counter[0] ),
    .B1(\simon0.tick_counter[2] ),
    .X(_0948_));
 sky130_fd_sc_hd__and3b_1 _3036_ (.A_N(_0947_),
    .B(_0948_),
    .C(_0943_),
    .X(_0949_));
 sky130_fd_sc_hd__clkbuf_1 _3037_ (.A(_0949_),
    .X(_0109_));
 sky130_fd_sc_hd__and2_1 _3038_ (.A(\simon0.tick_counter[3] ),
    .B(_0947_),
    .X(_0950_));
 sky130_fd_sc_hd__or2_1 _3039_ (.A(\simon0.tick_counter[3] ),
    .B(_0947_),
    .X(_0951_));
 sky130_fd_sc_hd__and3b_1 _3040_ (.A_N(_0950_),
    .B(_0951_),
    .C(_0943_),
    .X(_0952_));
 sky130_fd_sc_hd__clkbuf_1 _3041_ (.A(_0952_),
    .X(_0110_));
 sky130_fd_sc_hd__o21ai_1 _3042_ (.A1(\simon0.tick_counter[4] ),
    .A2(_0950_),
    .B1(_0944_),
    .Y(_0953_));
 sky130_fd_sc_hd__a21oi_1 _3043_ (.A1(\simon0.tick_counter[4] ),
    .A2(_0950_),
    .B1(_0953_),
    .Y(_0111_));
 sky130_fd_sc_hd__and3_1 _3044_ (.A(\simon0.tick_counter[4] ),
    .B(\simon0.tick_counter[5] ),
    .C(_0950_),
    .X(_0954_));
 sky130_fd_sc_hd__a31o_1 _3045_ (.A1(\simon0.tick_counter[3] ),
    .A2(\simon0.tick_counter[4] ),
    .A3(_0947_),
    .B1(\simon0.tick_counter[5] ),
    .X(_0955_));
 sky130_fd_sc_hd__and3b_1 _3046_ (.A_N(_0954_),
    .B(_0955_),
    .C(_0943_),
    .X(_0956_));
 sky130_fd_sc_hd__clkbuf_1 _3047_ (.A(_0956_),
    .X(_0112_));
 sky130_fd_sc_hd__and2_1 _3048_ (.A(\simon0.tick_counter[6] ),
    .B(_0954_),
    .X(_0957_));
 sky130_fd_sc_hd__o21ai_1 _3049_ (.A1(\simon0.tick_counter[6] ),
    .A2(_0954_),
    .B1(_0944_),
    .Y(_0958_));
 sky130_fd_sc_hd__nor2_1 _3050_ (.A(_0957_),
    .B(_0958_),
    .Y(_0113_));
 sky130_fd_sc_hd__and3_1 _3051_ (.A(\simon0.tick_counter[6] ),
    .B(\simon0.tick_counter[7] ),
    .C(_0954_),
    .X(_0959_));
 sky130_fd_sc_hd__o21ai_1 _3052_ (.A1(\simon0.tick_counter[7] ),
    .A2(_0957_),
    .B1(_0944_),
    .Y(_0960_));
 sky130_fd_sc_hd__nor2_1 _3053_ (.A(_0959_),
    .B(_0960_),
    .Y(_0114_));
 sky130_fd_sc_hd__and2_1 _3054_ (.A(\simon0.tick_counter[8] ),
    .B(_0959_),
    .X(_0961_));
 sky130_fd_sc_hd__inv_2 _3055_ (.A(_0961_),
    .Y(_0962_));
 sky130_fd_sc_hd__o211a_1 _3056_ (.A1(\simon0.tick_counter[8] ),
    .A2(_0959_),
    .B1(_0962_),
    .C1(_0944_),
    .X(_0115_));
 sky130_fd_sc_hd__and3_1 _3057_ (.A(\simon0.tick_counter[8] ),
    .B(\simon0.tick_counter[9] ),
    .C(_0959_),
    .X(_0963_));
 sky130_fd_sc_hd__o21ai_1 _3058_ (.A1(\simon0.tick_counter[9] ),
    .A2(_0961_),
    .B1(_0944_),
    .Y(_0964_));
 sky130_fd_sc_hd__nor2_1 _3059_ (.A(_0963_),
    .B(_0964_),
    .Y(_0116_));
 sky130_fd_sc_hd__o21ai_1 _3060_ (.A1(\simon0.tick_counter[10] ),
    .A2(_0963_),
    .B1(_0944_),
    .Y(_0965_));
 sky130_fd_sc_hd__a21oi_1 _3061_ (.A1(\simon0.tick_counter[10] ),
    .A2(_0963_),
    .B1(_0965_),
    .Y(_0117_));
 sky130_fd_sc_hd__and3_1 _3062_ (.A(\simon0.tick_counter[10] ),
    .B(\simon0.tick_counter[11] ),
    .C(_0963_),
    .X(_0966_));
 sky130_fd_sc_hd__a31o_1 _3063_ (.A1(\simon0.tick_counter[9] ),
    .A2(\simon0.tick_counter[10] ),
    .A3(_0961_),
    .B1(\simon0.tick_counter[11] ),
    .X(_0967_));
 sky130_fd_sc_hd__and3b_1 _3064_ (.A_N(_0966_),
    .B(_0943_),
    .C(_0967_),
    .X(_0968_));
 sky130_fd_sc_hd__clkbuf_1 _3065_ (.A(_0968_),
    .X(_0118_));
 sky130_fd_sc_hd__and2_1 _3066_ (.A(\simon0.tick_counter[12] ),
    .B(_0966_),
    .X(_0969_));
 sky130_fd_sc_hd__o21ai_1 _3067_ (.A1(\simon0.tick_counter[12] ),
    .A2(_0966_),
    .B1(_0944_),
    .Y(_0970_));
 sky130_fd_sc_hd__nor2_1 _3068_ (.A(_0969_),
    .B(_0970_),
    .Y(_0119_));
 sky130_fd_sc_hd__o21ai_1 _3069_ (.A1(\simon0.tick_counter[13] ),
    .A2(_0969_),
    .B1(_0944_),
    .Y(_0971_));
 sky130_fd_sc_hd__a21oi_1 _3070_ (.A1(\simon0.tick_counter[13] ),
    .A2(_0969_),
    .B1(_0971_),
    .Y(_0120_));
 sky130_fd_sc_hd__and3_1 _3071_ (.A(\simon0.tick_counter[13] ),
    .B(\simon0.tick_counter[14] ),
    .C(_0969_),
    .X(_0972_));
 sky130_fd_sc_hd__a31o_1 _3072_ (.A1(\simon0.tick_counter[12] ),
    .A2(\simon0.tick_counter[13] ),
    .A3(_0966_),
    .B1(\simon0.tick_counter[14] ),
    .X(_0973_));
 sky130_fd_sc_hd__and3b_1 _3073_ (.A_N(_0972_),
    .B(_0943_),
    .C(_0973_),
    .X(_0974_));
 sky130_fd_sc_hd__clkbuf_1 _3074_ (.A(_0974_),
    .X(_0121_));
 sky130_fd_sc_hd__a21boi_1 _3075_ (.A1(\simon0.tick_counter[15] ),
    .A2(_0972_),
    .B1_N(_0943_),
    .Y(_0975_));
 sky130_fd_sc_hd__o21a_1 _3076_ (.A1(\simon0.tick_counter[15] ),
    .A2(_0972_),
    .B1(_0975_),
    .X(_0122_));
 sky130_fd_sc_hd__a21bo_1 _3077_ (.A1(\simon0.state[4] ),
    .A2(_1170_),
    .B1_N(_1200_),
    .X(_0976_));
 sky130_fd_sc_hd__and2_1 _3078_ (.A(\simon0.seq_length[0] ),
    .B(_0976_),
    .X(_0977_));
 sky130_fd_sc_hd__nand2_1 _3079_ (.A(_1169_),
    .B(_0977_),
    .Y(_0978_));
 sky130_fd_sc_hd__o211a_1 _3080_ (.A1(\simon0.seq_length[0] ),
    .A2(_0976_),
    .B1(_0978_),
    .C1(_0499_),
    .X(_0123_));
 sky130_fd_sc_hd__or2_1 _3081_ (.A(\simon0.seq_length[1] ),
    .B(_0977_),
    .X(_0979_));
 sky130_fd_sc_hd__a21oi_2 _3082_ (.A1(\simon0.state[4] ),
    .A2(_1170_),
    .B1(net4),
    .Y(_0980_));
 sky130_fd_sc_hd__and3_1 _3083_ (.A(\simon0.seq_length[1] ),
    .B(\simon0.seq_length[0] ),
    .C(_0976_),
    .X(_0981_));
 sky130_fd_sc_hd__clkinv_2 _3084_ (.A(_0981_),
    .Y(_0982_));
 sky130_fd_sc_hd__and3_1 _3085_ (.A(_0979_),
    .B(_0980_),
    .C(_0982_),
    .X(_0983_));
 sky130_fd_sc_hd__clkbuf_1 _3086_ (.A(_0983_),
    .X(_0124_));
 sky130_fd_sc_hd__and2_1 _3087_ (.A(_1218_),
    .B(_0981_),
    .X(_0984_));
 sky130_fd_sc_hd__o21ai_1 _3088_ (.A1(_1218_),
    .A2(_0981_),
    .B1(_0980_),
    .Y(_0985_));
 sky130_fd_sc_hd__nor2_1 _3089_ (.A(_0984_),
    .B(_0985_),
    .Y(_0125_));
 sky130_fd_sc_hd__and3_1 _3090_ (.A(_1086_),
    .B(_1218_),
    .C(_0981_),
    .X(_0986_));
 sky130_fd_sc_hd__o21ai_1 _3091_ (.A1(_1086_),
    .A2(_0984_),
    .B1(_0980_),
    .Y(_0987_));
 sky130_fd_sc_hd__nor2_1 _3092_ (.A(_0986_),
    .B(_0987_),
    .Y(_0126_));
 sky130_fd_sc_hd__a21boi_1 _3093_ (.A1(_1217_),
    .A2(_0986_),
    .B1_N(_0980_),
    .Y(_0988_));
 sky130_fd_sc_hd__o21a_1 _3094_ (.A1(_1217_),
    .A2(_0986_),
    .B1(_0988_),
    .X(_0127_));
 sky130_fd_sc_hd__o21ba_1 _3095_ (.A1(\simon0.state[4] ),
    .A2(_1203_),
    .B1_N(_1189_),
    .X(_0989_));
 sky130_fd_sc_hd__o2111ai_4 _3096_ (.A1(_1170_),
    .A2(_1168_),
    .B1(_0834_),
    .C1(_1198_),
    .D1(_0989_),
    .Y(_0990_));
 sky130_fd_sc_hd__inv_2 _3097_ (.A(_0990_),
    .Y(_0991_));
 sky130_fd_sc_hd__o211ai_4 _3098_ (.A1(_1085_),
    .A2(_1169_),
    .B1(_1104_),
    .C1(_0991_),
    .Y(_0992_));
 sky130_fd_sc_hd__mux2_1 _3099_ (.A0(_0992_),
    .A1(_0991_),
    .S(\simon0.seq_counter[0] ),
    .X(_0993_));
 sky130_fd_sc_hd__nor2_1 _3100_ (.A(_1124_),
    .B(_0993_),
    .Y(_0128_));
 sky130_fd_sc_hd__o2bb2a_1 _3101_ (.A1_N(\simon0.seq_counter[1] ),
    .A2_N(_0990_),
    .B1(_0992_),
    .B2(_1098_),
    .X(_0994_));
 sky130_fd_sc_hd__nor2_1 _3102_ (.A(_1124_),
    .B(_0994_),
    .Y(_0129_));
 sky130_fd_sc_hd__o2bb2a_1 _3103_ (.A1_N(\simon0.seq_counter[2] ),
    .A2_N(_0990_),
    .B1(_0992_),
    .B2(_1095_),
    .X(_0995_));
 sky130_fd_sc_hd__nor2_1 _3104_ (.A(_1124_),
    .B(_0995_),
    .Y(_0130_));
 sky130_fd_sc_hd__o2bb2a_1 _3105_ (.A1_N(\simon0.seq_counter[3] ),
    .A2_N(_0990_),
    .B1(_0992_),
    .B2(_1090_),
    .X(_0996_));
 sky130_fd_sc_hd__nor2_1 _3106_ (.A(_1124_),
    .B(_0996_),
    .Y(_0131_));
 sky130_fd_sc_hd__nand2_1 _3107_ (.A(\simon0.seq_counter[4] ),
    .B(_0990_),
    .Y(_0997_));
 sky130_fd_sc_hd__or3b_1 _3108_ (.A(_1092_),
    .B(_0992_),
    .C_N(_1096_),
    .X(_0998_));
 sky130_fd_sc_hd__a21oi_1 _3109_ (.A1(_0997_),
    .A2(_0998_),
    .B1(_1201_),
    .Y(_0132_));
 sky130_fd_sc_hd__nor2_1 _3110_ (.A(_1169_),
    .B(\simon0.state[2] ),
    .Y(_0999_));
 sky130_fd_sc_hd__or2_1 _3111_ (.A(_1170_),
    .B(_0836_),
    .X(_1000_));
 sky130_fd_sc_hd__o21ai_2 _3112_ (.A1(_1169_),
    .A2(_0832_),
    .B1(_1000_),
    .Y(_1001_));
 sky130_fd_sc_hd__inv_2 _3113_ (.A(_1001_),
    .Y(_1002_));
 sky130_fd_sc_hd__or3_1 _3114_ (.A(\simon0.state[1] ),
    .B(\simon0.state[2] ),
    .C(_1205_),
    .X(_1003_));
 sky130_fd_sc_hd__o21ai_1 _3115_ (.A1(\simon0.millis_counter[8] ),
    .A2(\simon0.millis_counter[9] ),
    .B1(_1184_),
    .Y(_1004_));
 sky130_fd_sc_hd__nand2_1 _3116_ (.A(\simon0.millis_counter[7] ),
    .B(_1187_),
    .Y(_1005_));
 sky130_fd_sc_hd__o221a_1 _3117_ (.A1(_0999_),
    .A2(_1002_),
    .B1(_1003_),
    .B2(_1004_),
    .C1(_1005_),
    .X(_1006_));
 sky130_fd_sc_hd__clkinv_2 _3118_ (.A(\simon0.led[0] ),
    .Y(_1007_));
 sky130_fd_sc_hd__or2_2 _3119_ (.A(\simon0.state[4] ),
    .B(_0819_),
    .X(_1008_));
 sky130_fd_sc_hd__mux2_1 _3120_ (.A0(_1006_),
    .A1(_1007_),
    .S(_1008_),
    .X(_1009_));
 sky130_fd_sc_hd__nor2_1 _3121_ (.A(_1124_),
    .B(_1009_),
    .Y(_0133_));
 sky130_fd_sc_hd__mux2_1 _3122_ (.A0(_0833_),
    .A1(_0837_),
    .S(_1169_),
    .X(_1010_));
 sky130_fd_sc_hd__mux2_1 _3123_ (.A0(_1125_),
    .A1(_1147_),
    .S(_1170_),
    .X(_1011_));
 sky130_fd_sc_hd__and2_1 _3124_ (.A(_1005_),
    .B(_1003_),
    .X(_1012_));
 sky130_fd_sc_hd__o31a_1 _3125_ (.A1(_0999_),
    .A2(_1010_),
    .A3(_1011_),
    .B1(_1012_),
    .X(_1013_));
 sky130_fd_sc_hd__a21oi_1 _3126_ (.A1(_1109_),
    .A2(_1184_),
    .B1(_1003_),
    .Y(_1014_));
 sky130_fd_sc_hd__nand2_1 _3127_ (.A(\simon0.led[1] ),
    .B(_1008_),
    .Y(_1015_));
 sky130_fd_sc_hd__o31a_1 _3128_ (.A1(_1008_),
    .A2(_1013_),
    .A3(_1014_),
    .B1(_1015_),
    .X(_1016_));
 sky130_fd_sc_hd__nor2_1 _3129_ (.A(_1124_),
    .B(_1016_),
    .Y(_0134_));
 sky130_fd_sc_hd__or3b_1 _3130_ (.A(_0999_),
    .B(_1001_),
    .C_N(_1011_),
    .X(_1017_));
 sky130_fd_sc_hd__o21a_1 _3131_ (.A1(\simon0.millis_counter[8] ),
    .A2(_1108_),
    .B1(_1184_),
    .X(_1018_));
 sky130_fd_sc_hd__o2bb2a_1 _3132_ (.A1_N(_1012_),
    .A2_N(_1017_),
    .B1(_1018_),
    .B2(_1003_),
    .X(_1019_));
 sky130_fd_sc_hd__mux2_1 _3133_ (.A0(_1019_),
    .A1(\simon0.led[2] ),
    .S(_1008_),
    .X(_1020_));
 sky130_fd_sc_hd__and2_1 _3134_ (.A(_1084_),
    .B(_1020_),
    .X(_1021_));
 sky130_fd_sc_hd__clkbuf_1 _3135_ (.A(_1021_),
    .X(_0135_));
 sky130_fd_sc_hd__nand2_1 _3136_ (.A(\simon0.led[3] ),
    .B(_1008_),
    .Y(_1022_));
 sky130_fd_sc_hd__or3b_1 _3137_ (.A(_0999_),
    .B(_1001_),
    .C_N(_1010_),
    .X(_1023_));
 sky130_fd_sc_hd__a21oi_1 _3138_ (.A1(_1184_),
    .A2(_0803_),
    .B1(_1003_),
    .Y(_1024_));
 sky130_fd_sc_hd__a211o_1 _3139_ (.A1(_1012_),
    .A2(_1023_),
    .B1(_1024_),
    .C1(_1008_),
    .X(_1025_));
 sky130_fd_sc_hd__a21oi_1 _3140_ (.A1(_1022_),
    .A2(_1025_),
    .B1(_1201_),
    .Y(_0136_));
 sky130_fd_sc_hd__nand2_1 _3141_ (.A(_1252_),
    .B(_1244_),
    .Y(_1026_));
 sky130_fd_sc_hd__mux2_1 _3142_ (.A0(_1213_),
    .A1(\simon0.seq[30][0] ),
    .S(_1026_),
    .X(_1027_));
 sky130_fd_sc_hd__clkbuf_1 _3143_ (.A(_1027_),
    .X(_0137_));
 sky130_fd_sc_hd__mux2_1 _3144_ (.A0(_1223_),
    .A1(\simon0.seq[30][1] ),
    .S(_1026_),
    .X(_1028_));
 sky130_fd_sc_hd__clkbuf_1 _3145_ (.A(_1028_),
    .X(_0138_));
 sky130_fd_sc_hd__or2_1 _3146_ (.A(_1227_),
    .B(_1239_),
    .X(_1029_));
 sky130_fd_sc_hd__mux2_1 _3147_ (.A0(_1213_),
    .A1(\simon0.seq[19][0] ),
    .S(_1029_),
    .X(_1030_));
 sky130_fd_sc_hd__clkbuf_1 _3148_ (.A(_1030_),
    .X(_0139_));
 sky130_fd_sc_hd__mux2_1 _3149_ (.A0(_1223_),
    .A1(\simon0.seq[19][1] ),
    .S(_1029_),
    .X(_1031_));
 sky130_fd_sc_hd__clkbuf_1 _3150_ (.A(_1031_),
    .X(_0140_));
 sky130_fd_sc_hd__or3b_1 _3151_ (.A(_1218_),
    .B(_1225_),
    .C_N(_1217_),
    .X(_1032_));
 sky130_fd_sc_hd__or2_1 _3152_ (.A(_1278_),
    .B(_1032_),
    .X(_1033_));
 sky130_fd_sc_hd__mux2_1 _3153_ (.A0(_1231_),
    .A1(\simon0.seq[25][0] ),
    .S(_1033_),
    .X(_1034_));
 sky130_fd_sc_hd__clkbuf_1 _3154_ (.A(_1034_),
    .X(_0141_));
 sky130_fd_sc_hd__mux2_1 _3155_ (.A0(_1236_),
    .A1(\simon0.seq[25][1] ),
    .S(_1033_),
    .X(_1035_));
 sky130_fd_sc_hd__clkbuf_1 _3156_ (.A(_1035_),
    .X(_0142_));
 sky130_fd_sc_hd__nor2_1 _3157_ (.A(_1238_),
    .B(_1032_),
    .Y(_1036_));
 sky130_fd_sc_hd__mux2_1 _3158_ (.A0(\simon0.seq[24][0] ),
    .A1(_1273_),
    .S(_1036_),
    .X(_1037_));
 sky130_fd_sc_hd__clkbuf_1 _3159_ (.A(_1037_),
    .X(_0143_));
 sky130_fd_sc_hd__mux2_1 _3160_ (.A0(\simon0.seq[24][1] ),
    .A1(_1276_),
    .S(_1036_),
    .X(_1038_));
 sky130_fd_sc_hd__clkbuf_1 _3161_ (.A(_1038_),
    .X(_0144_));
 sky130_fd_sc_hd__nand2_1 _3162_ (.A(_1248_),
    .B(_1289_),
    .Y(_1039_));
 sky130_fd_sc_hd__mux2_1 _3163_ (.A0(_1231_),
    .A1(\simon0.seq[23][0] ),
    .S(_1039_),
    .X(_1040_));
 sky130_fd_sc_hd__clkbuf_1 _3164_ (.A(_1040_),
    .X(_0145_));
 sky130_fd_sc_hd__mux2_1 _3165_ (.A0(_1236_),
    .A1(\simon0.seq[23][1] ),
    .S(_1039_),
    .X(_1041_));
 sky130_fd_sc_hd__clkbuf_1 _3166_ (.A(_1041_),
    .X(_0146_));
 sky130_fd_sc_hd__nor2_1 _3167_ (.A(_1233_),
    .B(_1032_),
    .Y(_1042_));
 sky130_fd_sc_hd__mux2_1 _3168_ (.A0(\simon0.seq[26][0] ),
    .A1(_1273_),
    .S(_1042_),
    .X(_1043_));
 sky130_fd_sc_hd__clkbuf_1 _3169_ (.A(_1043_),
    .X(_0147_));
 sky130_fd_sc_hd__mux2_1 _3170_ (.A0(\simon0.seq[26][1] ),
    .A1(_1276_),
    .S(_1042_),
    .X(_1044_));
 sky130_fd_sc_hd__clkbuf_1 _3171_ (.A(_1044_),
    .X(_0148_));
 sky130_fd_sc_hd__nand2_1 _3172_ (.A(_1216_),
    .B(_1244_),
    .Y(_1045_));
 sky130_fd_sc_hd__mux2_1 _3173_ (.A0(_1231_),
    .A1(\simon0.seq[28][0] ),
    .S(_1045_),
    .X(_1046_));
 sky130_fd_sc_hd__clkbuf_1 _3174_ (.A(_1046_),
    .X(_0149_));
 sky130_fd_sc_hd__mux2_1 _3175_ (.A0(_1236_),
    .A1(\simon0.seq[28][1] ),
    .S(_1045_),
    .X(_1047_));
 sky130_fd_sc_hd__clkbuf_1 _3176_ (.A(_1047_),
    .X(_0150_));
 sky130_fd_sc_hd__nor2_1 _3177_ (.A(_1278_),
    .B(_1285_),
    .Y(_1048_));
 sky130_fd_sc_hd__mux2_1 _3178_ (.A0(\simon0.seq[1][0] ),
    .A1(_1273_),
    .S(_1048_),
    .X(_1049_));
 sky130_fd_sc_hd__clkbuf_1 _3179_ (.A(_1049_),
    .X(_0151_));
 sky130_fd_sc_hd__mux2_1 _3180_ (.A0(\simon0.seq[1][1] ),
    .A1(_1276_),
    .S(_1048_),
    .X(_1050_));
 sky130_fd_sc_hd__clkbuf_1 _3181_ (.A(_1050_),
    .X(_0152_));
 sky130_fd_sc_hd__nor2_1 _3182_ (.A(_1265_),
    .B(_1032_),
    .Y(_1051_));
 sky130_fd_sc_hd__mux2_1 _3183_ (.A0(\simon0.seq[27][0] ),
    .A1(_1273_),
    .S(_1051_),
    .X(_1052_));
 sky130_fd_sc_hd__clkbuf_1 _3184_ (.A(_1052_),
    .X(_0153_));
 sky130_fd_sc_hd__mux2_1 _3185_ (.A0(\simon0.seq[27][1] ),
    .A1(_1276_),
    .S(_1051_),
    .X(_1053_));
 sky130_fd_sc_hd__clkbuf_1 _3186_ (.A(_1053_),
    .X(_0154_));
 sky130_fd_sc_hd__nor2_1 _3187_ (.A(_1233_),
    .B(_1285_),
    .Y(_1054_));
 sky130_fd_sc_hd__mux2_1 _3188_ (.A0(\simon0.seq[2][0] ),
    .A1(_1273_),
    .S(_1054_),
    .X(_1055_));
 sky130_fd_sc_hd__clkbuf_1 _3189_ (.A(_1055_),
    .X(_0155_));
 sky130_fd_sc_hd__mux2_1 _3190_ (.A0(\simon0.seq[2][1] ),
    .A1(_1276_),
    .S(_1054_),
    .X(_1056_));
 sky130_fd_sc_hd__clkbuf_1 _3191_ (.A(_1056_),
    .X(_0156_));
 sky130_fd_sc_hd__nor2_1 _3192_ (.A(_1226_),
    .B(_1278_),
    .Y(_1057_));
 sky130_fd_sc_hd__mux2_1 _3193_ (.A0(\simon0.seq[9][0] ),
    .A1(_1273_),
    .S(_1057_),
    .X(_1058_));
 sky130_fd_sc_hd__clkbuf_1 _3194_ (.A(_1058_),
    .X(_0157_));
 sky130_fd_sc_hd__mux2_1 _3195_ (.A0(\simon0.seq[9][1] ),
    .A1(_1276_),
    .S(_1057_),
    .X(_1059_));
 sky130_fd_sc_hd__clkbuf_1 _3196_ (.A(_1059_),
    .X(_0158_));
 sky130_fd_sc_hd__nor2_1 _3197_ (.A(_1233_),
    .B(_1239_),
    .Y(_1060_));
 sky130_fd_sc_hd__mux2_1 _3198_ (.A0(\simon0.seq[18][0] ),
    .A1(_1212_),
    .S(_1060_),
    .X(_1061_));
 sky130_fd_sc_hd__clkbuf_1 _3199_ (.A(_1061_),
    .X(_0159_));
 sky130_fd_sc_hd__mux2_1 _3200_ (.A0(\simon0.seq[18][1] ),
    .A1(_1222_),
    .S(_1060_),
    .X(_1062_));
 sky130_fd_sc_hd__clkbuf_1 _3201_ (.A(_1062_),
    .X(_0160_));
 sky130_fd_sc_hd__nand2_1 _3202_ (.A(_1248_),
    .B(_1244_),
    .Y(_1063_));
 sky130_fd_sc_hd__mux2_1 _3203_ (.A0(_1231_),
    .A1(\simon0.seq[31][0] ),
    .S(_1063_),
    .X(_1064_));
 sky130_fd_sc_hd__clkbuf_1 _3204_ (.A(_1064_),
    .X(_0161_));
 sky130_fd_sc_hd__mux2_1 _3205_ (.A0(_1236_),
    .A1(\simon0.seq[31][1] ),
    .S(_1063_),
    .X(_1065_));
 sky130_fd_sc_hd__clkbuf_1 _3206_ (.A(_1065_),
    .X(_0162_));
 sky130_fd_sc_hd__nor2_1 _3207_ (.A(_1201_),
    .B(_0993_),
    .Y(_0163_));
 sky130_fd_sc_hd__nor2_1 _3208_ (.A(_1201_),
    .B(_0994_),
    .Y(_0164_));
 sky130_fd_sc_hd__nor2_1 _3209_ (.A(_1201_),
    .B(_0995_),
    .Y(_0165_));
 sky130_fd_sc_hd__nor2_1 _3210_ (.A(_1201_),
    .B(_0996_),
    .Y(_0166_));
 sky130_fd_sc_hd__a21oi_1 _3211_ (.A1(_0997_),
    .A2(_0998_),
    .B1(_1201_),
    .Y(_0167_));
 sky130_fd_sc_hd__nand2_1 _3212_ (.A(_1243_),
    .B(_1289_),
    .Y(_1066_));
 sky130_fd_sc_hd__mux2_1 _3213_ (.A0(_1231_),
    .A1(\simon0.seq[21][0] ),
    .S(_1066_),
    .X(_1067_));
 sky130_fd_sc_hd__clkbuf_1 _3214_ (.A(_1067_),
    .X(_0168_));
 sky130_fd_sc_hd__mux2_1 _3215_ (.A0(_1236_),
    .A1(\simon0.seq[21][1] ),
    .S(_1066_),
    .X(_1068_));
 sky130_fd_sc_hd__clkbuf_1 _3216_ (.A(_1068_),
    .X(_0169_));
 sky130_fd_sc_hd__nor2_1 _3217_ (.A(_1239_),
    .B(_1278_),
    .Y(_1069_));
 sky130_fd_sc_hd__mux2_1 _3218_ (.A0(\simon0.seq[17][0] ),
    .A1(_1212_),
    .S(_1069_),
    .X(_1070_));
 sky130_fd_sc_hd__clkbuf_1 _3219_ (.A(_1070_),
    .X(_0170_));
 sky130_fd_sc_hd__mux2_1 _3220_ (.A0(\simon0.seq[17][1] ),
    .A1(_1222_),
    .S(_1069_),
    .X(_1071_));
 sky130_fd_sc_hd__clkbuf_1 _3221_ (.A(_1071_),
    .X(_0171_));
 sky130_fd_sc_hd__dfxtp_1 _3222_ (.CLK(clknet_4_7_0_wb_clk_i),
    .D(_0013_),
    .Q(\simon0.seq[12][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3223_ (.CLK(clknet_4_6_0_wb_clk_i),
    .D(_0014_),
    .Q(\simon0.seq[12][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3224_ (.CLK(clknet_4_5_0_wb_clk_i),
    .D(_0015_),
    .Q(\simon0.seq[11][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3225_ (.CLK(clknet_4_5_0_wb_clk_i),
    .D(_0016_),
    .Q(\simon0.seq[11][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3226_ (.CLK(clknet_4_5_0_wb_clk_i),
    .D(_0017_),
    .Q(\simon0.seq[10][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3227_ (.CLK(clknet_4_5_0_wb_clk_i),
    .D(_0018_),
    .Q(\simon0.seq[10][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3228_ (.CLK(clknet_4_3_0_wb_clk_i),
    .D(_0019_),
    .Q(\simon0.seq[16][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3229_ (.CLK(clknet_4_3_0_wb_clk_i),
    .D(_0020_),
    .Q(\simon0.seq[16][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3230_ (.CLK(clknet_4_7_0_wb_clk_i),
    .D(_0021_),
    .Q(\simon0.seq[29][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3231_ (.CLK(clknet_4_7_0_wb_clk_i),
    .D(_0022_),
    .Q(\simon0.seq[29][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3232_ (.CLK(clknet_4_7_0_wb_clk_i),
    .D(_0023_),
    .Q(\simon0.seq[15][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3233_ (.CLK(clknet_4_7_0_wb_clk_i),
    .D(_0024_),
    .Q(\simon0.seq[15][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3234_ (.CLK(clknet_4_7_0_wb_clk_i),
    .D(_0025_),
    .Q(\simon0.seq[14][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3235_ (.CLK(clknet_4_7_0_wb_clk_i),
    .D(_0026_),
    .Q(\simon0.seq[14][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3236_ (.CLK(clknet_4_7_0_wb_clk_i),
    .D(_0027_),
    .Q(\simon0.seq[13][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3237_ (.CLK(clknet_4_6_0_wb_clk_i),
    .D(_0028_),
    .Q(\simon0.seq[13][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3238_ (.CLK(clknet_4_5_0_wb_clk_i),
    .D(_0029_),
    .Q(\simon0.seq[8][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3239_ (.CLK(clknet_4_5_0_wb_clk_i),
    .D(_0030_),
    .Q(\simon0.seq[8][1] ));
 sky130_fd_sc_hd__dfxtp_2 _3240_ (.CLK(clknet_4_13_0_wb_clk_i),
    .D(_0031_),
    .Q(\simon0.user_input[0] ));
 sky130_fd_sc_hd__dfxtp_1 _3241_ (.CLK(clknet_4_13_0_wb_clk_i),
    .D(_0032_),
    .Q(\simon0.user_input[1] ));
 sky130_fd_sc_hd__dfxtp_1 _3242_ (.CLK(clknet_4_4_0_wb_clk_i),
    .D(_0033_),
    .Q(\simon0.seq[7][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3243_ (.CLK(clknet_4_1_0_wb_clk_i),
    .D(_0034_),
    .Q(\simon0.seq[7][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3244_ (.CLK(clknet_4_5_0_wb_clk_i),
    .D(_0035_),
    .Q(\simon0.seq[6][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3245_ (.CLK(clknet_4_5_0_wb_clk_i),
    .D(_0036_),
    .Q(\simon0.seq[6][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3246_ (.CLK(clknet_4_13_0_wb_clk_i),
    .D(_0005_),
    .Q(\simon0.state[0] ));
 sky130_fd_sc_hd__dfxtp_1 _3247_ (.CLK(clknet_4_13_0_wb_clk_i),
    .D(_0006_),
    .Q(\simon0.state[1] ));
 sky130_fd_sc_hd__dfxtp_1 _3248_ (.CLK(clknet_4_13_0_wb_clk_i),
    .D(_0007_),
    .Q(\simon0.state[2] ));
 sky130_fd_sc_hd__dfxtp_1 _3249_ (.CLK(clknet_4_13_0_wb_clk_i),
    .D(_0008_),
    .Q(\simon0.state[3] ));
 sky130_fd_sc_hd__dfxtp_2 _3250_ (.CLK(clknet_4_13_0_wb_clk_i),
    .D(_0009_),
    .Q(\simon0.state[4] ));
 sky130_fd_sc_hd__dfxtp_1 _3251_ (.CLK(clknet_4_13_0_wb_clk_i),
    .D(_0010_),
    .Q(\simon0.state[5] ));
 sky130_fd_sc_hd__dfxtp_1 _3252_ (.CLK(clknet_4_13_0_wb_clk_i),
    .D(_0011_),
    .Q(\simon0.state[6] ));
 sky130_fd_sc_hd__dfxtp_2 _3253_ (.CLK(clknet_4_6_0_wb_clk_i),
    .D(_0012_),
    .Q(\simon0.state[7] ));
 sky130_fd_sc_hd__dfxtp_1 _3254_ (.CLK(clknet_4_3_0_wb_clk_i),
    .D(_0037_),
    .Q(\simon0.seq[0][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3255_ (.CLK(clknet_4_0_0_wb_clk_i),
    .D(_0038_),
    .Q(\simon0.seq[0][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3256_ (.CLK(clknet_4_4_0_wb_clk_i),
    .D(_0039_),
    .Q(\simon0.seq[5][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3257_ (.CLK(clknet_4_1_0_wb_clk_i),
    .D(_0040_),
    .Q(\simon0.seq[5][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3258_ (.CLK(clknet_4_4_0_wb_clk_i),
    .D(_0041_),
    .Q(\simon0.seq[4][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3259_ (.CLK(clknet_4_1_0_wb_clk_i),
    .D(_0042_),
    .Q(\simon0.seq[4][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3260_ (.CLK(clknet_4_1_0_wb_clk_i),
    .D(_0043_),
    .Q(\simon0.seq[3][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3261_ (.CLK(clknet_4_0_0_wb_clk_i),
    .D(_0044_),
    .Q(\simon0.seq[3][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3262_ (.CLK(clknet_4_4_0_wb_clk_i),
    .D(_0045_),
    .Q(\simon0.seq[22][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3263_ (.CLK(clknet_4_4_0_wb_clk_i),
    .D(_0046_),
    .Q(\simon0.seq[22][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3264_ (.CLK(clknet_4_12_0_wb_clk_i),
    .D(_0047_),
    .Q(\simon0.play1.tick_counter[0] ));
 sky130_fd_sc_hd__dfxtp_1 _3265_ (.CLK(clknet_4_12_0_wb_clk_i),
    .D(_0048_),
    .Q(\simon0.play1.tick_counter[1] ));
 sky130_fd_sc_hd__dfxtp_1 _3266_ (.CLK(clknet_4_9_0_wb_clk_i),
    .D(_0049_),
    .Q(\simon0.play1.tick_counter[2] ));
 sky130_fd_sc_hd__dfxtp_1 _3267_ (.CLK(clknet_4_9_0_wb_clk_i),
    .D(_0050_),
    .Q(\simon0.play1.tick_counter[3] ));
 sky130_fd_sc_hd__dfxtp_1 _3268_ (.CLK(clknet_4_9_0_wb_clk_i),
    .D(_0051_),
    .Q(\simon0.play1.tick_counter[4] ));
 sky130_fd_sc_hd__dfxtp_1 _3269_ (.CLK(clknet_4_9_0_wb_clk_i),
    .D(_0052_),
    .Q(\simon0.play1.tick_counter[5] ));
 sky130_fd_sc_hd__dfxtp_1 _3270_ (.CLK(clknet_4_9_0_wb_clk_i),
    .D(_0053_),
    .Q(\simon0.play1.tick_counter[6] ));
 sky130_fd_sc_hd__dfxtp_1 _3271_ (.CLK(clknet_4_11_0_wb_clk_i),
    .D(_0054_),
    .Q(\simon0.play1.tick_counter[7] ));
 sky130_fd_sc_hd__dfxtp_1 _3272_ (.CLK(clknet_4_11_0_wb_clk_i),
    .D(_0055_),
    .Q(\simon0.play1.tick_counter[8] ));
 sky130_fd_sc_hd__dfxtp_1 _3273_ (.CLK(clknet_4_9_0_wb_clk_i),
    .D(_0056_),
    .Q(\simon0.play1.tick_counter[9] ));
 sky130_fd_sc_hd__dfxtp_1 _3274_ (.CLK(clknet_4_8_0_wb_clk_i),
    .D(_0057_),
    .Q(\simon0.play1.tick_counter[10] ));
 sky130_fd_sc_hd__dfxtp_1 _3275_ (.CLK(clknet_4_8_0_wb_clk_i),
    .D(_0058_),
    .Q(\simon0.play1.tick_counter[11] ));
 sky130_fd_sc_hd__dfxtp_1 _3276_ (.CLK(clknet_4_2_0_wb_clk_i),
    .D(_0059_),
    .Q(\simon0.play1.tick_counter[12] ));
 sky130_fd_sc_hd__dfxtp_1 _3277_ (.CLK(clknet_4_8_0_wb_clk_i),
    .D(_0060_),
    .Q(\simon0.play1.tick_counter[13] ));
 sky130_fd_sc_hd__dfxtp_1 _3278_ (.CLK(clknet_4_8_0_wb_clk_i),
    .D(_0061_),
    .Q(\simon0.play1.tick_counter[14] ));
 sky130_fd_sc_hd__dfxtp_1 _3279_ (.CLK(clknet_4_8_0_wb_clk_i),
    .D(_0062_),
    .Q(\simon0.play1.tick_counter[15] ));
 sky130_fd_sc_hd__dfxtp_1 _3280_ (.CLK(clknet_4_8_0_wb_clk_i),
    .D(_0063_),
    .Q(\simon0.play1.tick_counter[16] ));
 sky130_fd_sc_hd__dfxtp_1 _3281_ (.CLK(clknet_4_8_0_wb_clk_i),
    .D(_0064_),
    .Q(\simon0.play1.tick_counter[17] ));
 sky130_fd_sc_hd__dfxtp_1 _3282_ (.CLK(clknet_4_8_0_wb_clk_i),
    .D(_0065_),
    .Q(\simon0.play1.tick_counter[18] ));
 sky130_fd_sc_hd__dfxtp_1 _3283_ (.CLK(clknet_4_10_0_wb_clk_i),
    .D(_0066_),
    .Q(\simon0.play1.tick_counter[19] ));
 sky130_fd_sc_hd__dfxtp_1 _3284_ (.CLK(clknet_4_10_0_wb_clk_i),
    .D(_0067_),
    .Q(\simon0.play1.tick_counter[20] ));
 sky130_fd_sc_hd__dfxtp_2 _3285_ (.CLK(clknet_4_10_0_wb_clk_i),
    .D(_0068_),
    .Q(\simon0.play1.tick_counter[21] ));
 sky130_fd_sc_hd__dfxtp_1 _3286_ (.CLK(clknet_4_10_0_wb_clk_i),
    .D(_0069_),
    .Q(\simon0.play1.tick_counter[22] ));
 sky130_fd_sc_hd__dfxtp_1 _3287_ (.CLK(clknet_4_10_0_wb_clk_i),
    .D(_0070_),
    .Q(\simon0.play1.tick_counter[23] ));
 sky130_fd_sc_hd__dfxtp_1 _3288_ (.CLK(clknet_4_10_0_wb_clk_i),
    .D(_0071_),
    .Q(\simon0.play1.tick_counter[24] ));
 sky130_fd_sc_hd__dfxtp_1 _3289_ (.CLK(clknet_4_10_0_wb_clk_i),
    .D(_0072_),
    .Q(\simon0.play1.tick_counter[25] ));
 sky130_fd_sc_hd__dfxtp_1 _3290_ (.CLK(clknet_4_10_0_wb_clk_i),
    .D(_0073_),
    .Q(\simon0.play1.tick_counter[26] ));
 sky130_fd_sc_hd__dfxtp_1 _3291_ (.CLK(clknet_4_10_0_wb_clk_i),
    .D(_0074_),
    .Q(\simon0.play1.tick_counter[27] ));
 sky130_fd_sc_hd__dfxtp_1 _3292_ (.CLK(clknet_4_11_0_wb_clk_i),
    .D(_0075_),
    .Q(\simon0.play1.tick_counter[28] ));
 sky130_fd_sc_hd__dfxtp_1 _3293_ (.CLK(clknet_4_11_0_wb_clk_i),
    .D(_0076_),
    .Q(\simon0.play1.tick_counter[29] ));
 sky130_fd_sc_hd__dfxtp_1 _3294_ (.CLK(clknet_4_11_0_wb_clk_i),
    .D(_0077_),
    .Q(\simon0.play1.tick_counter[30] ));
 sky130_fd_sc_hd__dfxtp_1 _3295_ (.CLK(clknet_4_10_0_wb_clk_i),
    .D(_0078_),
    .Q(\simon0.play1.tick_counter[31] ));
 sky130_fd_sc_hd__dfxtp_1 _3296_ (.CLK(clknet_4_11_0_wb_clk_i),
    .D(_0079_),
    .Q(\simon0.play1.sound ));
 sky130_fd_sc_hd__dfxtp_1 _3297_ (.CLK(clknet_4_6_0_wb_clk_i),
    .D(_0080_),
    .Q(\simon0.seq[20][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3298_ (.CLK(clknet_4_6_0_wb_clk_i),
    .D(_0081_),
    .Q(\simon0.seq[20][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3299_ (.CLK(clknet_4_6_0_wb_clk_i),
    .D(_0082_),
    .Q(\simon0.next_random[0] ));
 sky130_fd_sc_hd__dfxtp_1 _3300_ (.CLK(clknet_4_6_0_wb_clk_i),
    .D(_0083_),
    .Q(\simon0.next_random[1] ));
 sky130_fd_sc_hd__dfxtp_2 _3301_ (.CLK(clknet_4_14_0_wb_clk_i),
    .D(_0084_),
    .Q(\simon0.tone_sequence_counter[0] ));
 sky130_fd_sc_hd__dfxtp_2 _3302_ (.CLK(clknet_4_14_0_wb_clk_i),
    .D(_0085_),
    .Q(\simon0.tone_sequence_counter[1] ));
 sky130_fd_sc_hd__dfxtp_1 _3303_ (.CLK(clknet_4_14_0_wb_clk_i),
    .D(_0086_),
    .Q(\simon0.tone_sequence_counter[2] ));
 sky130_fd_sc_hd__dfxtp_1 _3304_ (.CLK(clknet_4_12_0_wb_clk_i),
    .D(_0087_),
    .Q(\simon0.play1.freq[0] ));
 sky130_fd_sc_hd__dfxtp_1 _3305_ (.CLK(clknet_4_12_0_wb_clk_i),
    .D(_0088_),
    .Q(\simon0.play1.freq[1] ));
 sky130_fd_sc_hd__dfxtp_1 _3306_ (.CLK(clknet_4_12_0_wb_clk_i),
    .D(_0089_),
    .Q(\simon0.play1.freq[2] ));
 sky130_fd_sc_hd__dfxtp_1 _3307_ (.CLK(clknet_4_12_0_wb_clk_i),
    .D(_0090_),
    .Q(\simon0.play1.freq[3] ));
 sky130_fd_sc_hd__dfxtp_1 _3308_ (.CLK(clknet_4_14_0_wb_clk_i),
    .D(_0091_),
    .Q(\simon0.play1.freq[4] ));
 sky130_fd_sc_hd__dfxtp_1 _3309_ (.CLK(clknet_4_11_0_wb_clk_i),
    .D(_0092_),
    .Q(\simon0.play1.freq[5] ));
 sky130_fd_sc_hd__dfxtp_1 _3310_ (.CLK(clknet_4_9_0_wb_clk_i),
    .D(_0093_),
    .Q(\simon0.play1.freq[6] ));
 sky130_fd_sc_hd__dfxtp_1 _3311_ (.CLK(clknet_4_12_0_wb_clk_i),
    .D(_0094_),
    .Q(\simon0.play1.freq[7] ));
 sky130_fd_sc_hd__dfxtp_2 _3312_ (.CLK(clknet_4_12_0_wb_clk_i),
    .D(_0095_),
    .Q(\simon0.play1.freq[8] ));
 sky130_fd_sc_hd__dfxtp_2 _3313_ (.CLK(clknet_4_14_0_wb_clk_i),
    .D(_0096_),
    .Q(\simon0.play1.freq[9] ));
 sky130_fd_sc_hd__dfxtp_1 _3314_ (.CLK(clknet_4_14_0_wb_clk_i),
    .D(_0097_),
    .Q(\simon0.millis_counter[0] ));
 sky130_fd_sc_hd__dfxtp_1 _3315_ (.CLK(clknet_4_14_0_wb_clk_i),
    .D(_0098_),
    .Q(\simon0.millis_counter[1] ));
 sky130_fd_sc_hd__dfxtp_1 _3316_ (.CLK(clknet_4_15_0_wb_clk_i),
    .D(_0099_),
    .Q(\simon0.millis_counter[2] ));
 sky130_fd_sc_hd__dfxtp_1 _3317_ (.CLK(clknet_4_15_0_wb_clk_i),
    .D(_0100_),
    .Q(\simon0.millis_counter[3] ));
 sky130_fd_sc_hd__dfxtp_2 _3318_ (.CLK(clknet_4_15_0_wb_clk_i),
    .D(_0101_),
    .Q(\simon0.millis_counter[4] ));
 sky130_fd_sc_hd__dfxtp_1 _3319_ (.CLK(clknet_4_15_0_wb_clk_i),
    .D(_0102_),
    .Q(\simon0.millis_counter[5] ));
 sky130_fd_sc_hd__dfxtp_1 _3320_ (.CLK(clknet_4_15_0_wb_clk_i),
    .D(_0103_),
    .Q(\simon0.millis_counter[6] ));
 sky130_fd_sc_hd__dfxtp_1 _3321_ (.CLK(clknet_4_15_0_wb_clk_i),
    .D(_0104_),
    .Q(\simon0.millis_counter[7] ));
 sky130_fd_sc_hd__dfxtp_1 _3322_ (.CLK(clknet_4_15_0_wb_clk_i),
    .D(_0105_),
    .Q(\simon0.millis_counter[8] ));
 sky130_fd_sc_hd__dfxtp_1 _3323_ (.CLK(clknet_4_15_0_wb_clk_i),
    .D(_0106_),
    .Q(\simon0.millis_counter[9] ));
 sky130_fd_sc_hd__dfxtp_1 _3324_ (.CLK(clknet_4_2_0_wb_clk_i),
    .D(_0107_),
    .Q(\simon0.tick_counter[0] ));
 sky130_fd_sc_hd__dfxtp_1 _3325_ (.CLK(clknet_4_2_0_wb_clk_i),
    .D(_0108_),
    .Q(\simon0.tick_counter[1] ));
 sky130_fd_sc_hd__dfxtp_1 _3326_ (.CLK(clknet_4_2_0_wb_clk_i),
    .D(_0109_),
    .Q(\simon0.tick_counter[2] ));
 sky130_fd_sc_hd__dfxtp_1 _3327_ (.CLK(clknet_4_0_0_wb_clk_i),
    .D(_0110_),
    .Q(\simon0.tick_counter[3] ));
 sky130_fd_sc_hd__dfxtp_1 _3328_ (.CLK(clknet_4_0_0_wb_clk_i),
    .D(_0111_),
    .Q(\simon0.tick_counter[4] ));
 sky130_fd_sc_hd__dfxtp_1 _3329_ (.CLK(clknet_4_0_0_wb_clk_i),
    .D(_0112_),
    .Q(\simon0.tick_counter[5] ));
 sky130_fd_sc_hd__dfxtp_1 _3330_ (.CLK(clknet_4_0_0_wb_clk_i),
    .D(_0113_),
    .Q(\simon0.tick_counter[6] ));
 sky130_fd_sc_hd__dfxtp_1 _3331_ (.CLK(clknet_4_0_0_wb_clk_i),
    .D(_0114_),
    .Q(\simon0.tick_counter[7] ));
 sky130_fd_sc_hd__dfxtp_1 _3332_ (.CLK(clknet_4_0_0_wb_clk_i),
    .D(_0115_),
    .Q(\simon0.tick_counter[8] ));
 sky130_fd_sc_hd__dfxtp_1 _3333_ (.CLK(clknet_4_0_0_wb_clk_i),
    .D(_0116_),
    .Q(\simon0.tick_counter[9] ));
 sky130_fd_sc_hd__dfxtp_1 _3334_ (.CLK(clknet_4_0_0_wb_clk_i),
    .D(_0117_),
    .Q(\simon0.tick_counter[10] ));
 sky130_fd_sc_hd__dfxtp_1 _3335_ (.CLK(clknet_4_0_0_wb_clk_i),
    .D(_0118_),
    .Q(\simon0.tick_counter[11] ));
 sky130_fd_sc_hd__dfxtp_1 _3336_ (.CLK(clknet_4_0_0_wb_clk_i),
    .D(_0119_),
    .Q(\simon0.tick_counter[12] ));
 sky130_fd_sc_hd__dfxtp_1 _3337_ (.CLK(clknet_4_0_0_wb_clk_i),
    .D(_0120_),
    .Q(\simon0.tick_counter[13] ));
 sky130_fd_sc_hd__dfxtp_1 _3338_ (.CLK(clknet_4_2_0_wb_clk_i),
    .D(_0121_),
    .Q(\simon0.tick_counter[14] ));
 sky130_fd_sc_hd__dfxtp_1 _3339_ (.CLK(clknet_4_2_0_wb_clk_i),
    .D(_0122_),
    .Q(\simon0.tick_counter[15] ));
 sky130_fd_sc_hd__dfxtp_2 _3340_ (.CLK(clknet_4_6_0_wb_clk_i),
    .D(_0123_),
    .Q(\simon0.seq_length[0] ));
 sky130_fd_sc_hd__dfxtp_2 _3341_ (.CLK(clknet_4_6_0_wb_clk_i),
    .D(_0124_),
    .Q(\simon0.seq_length[1] ));
 sky130_fd_sc_hd__dfxtp_1 _3342_ (.CLK(clknet_4_3_0_wb_clk_i),
    .D(_0125_),
    .Q(\simon0.seq_length[2] ));
 sky130_fd_sc_hd__dfxtp_1 _3343_ (.CLK(clknet_4_3_0_wb_clk_i),
    .D(_0126_),
    .Q(\simon0.seq_length[3] ));
 sky130_fd_sc_hd__dfxtp_1 _3344_ (.CLK(clknet_4_3_0_wb_clk_i),
    .D(_0127_),
    .Q(\simon0.seq_length[4] ));
 sky130_fd_sc_hd__dfxtp_1 _3345_ (.CLK(clknet_4_6_0_wb_clk_i),
    .D(_0128_),
    .Q(\simon0.seq_counter[0] ));
 sky130_fd_sc_hd__dfxtp_1 _3346_ (.CLK(clknet_4_3_0_wb_clk_i),
    .D(_0129_),
    .Q(\simon0.seq_counter[1] ));
 sky130_fd_sc_hd__dfxtp_1 _3347_ (.CLK(clknet_4_3_0_wb_clk_i),
    .D(_0130_),
    .Q(\simon0.seq_counter[2] ));
 sky130_fd_sc_hd__dfxtp_1 _3348_ (.CLK(clknet_4_6_0_wb_clk_i),
    .D(_0131_),
    .Q(\simon0.seq_counter[3] ));
 sky130_fd_sc_hd__dfxtp_1 _3349_ (.CLK(clknet_4_2_0_wb_clk_i),
    .D(_0132_),
    .Q(\simon0.seq_counter[4] ));
 sky130_fd_sc_hd__dfxtp_4 _3350_ (.CLK(clknet_4_13_0_wb_clk_i),
    .D(_0133_),
    .Q(\simon0.led[0] ));
 sky130_fd_sc_hd__dfxtp_2 _3351_ (.CLK(clknet_4_13_0_wb_clk_i),
    .D(_0134_),
    .Q(\simon0.led[1] ));
 sky130_fd_sc_hd__dfxtp_1 _3352_ (.CLK(clknet_4_15_0_wb_clk_i),
    .D(_0135_),
    .Q(\simon0.led[2] ));
 sky130_fd_sc_hd__dfxtp_1 _3353_ (.CLK(clknet_4_13_0_wb_clk_i),
    .D(_0136_),
    .Q(\simon0.led[3] ));
 sky130_fd_sc_hd__dfxtp_1 _3354_ (.CLK(clknet_4_5_0_wb_clk_i),
    .D(_0137_),
    .Q(\simon0.seq[30][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3355_ (.CLK(clknet_4_5_0_wb_clk_i),
    .D(_0138_),
    .Q(\simon0.seq[30][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3356_ (.CLK(clknet_4_3_0_wb_clk_i),
    .D(_0139_),
    .Q(\simon0.seq[19][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3357_ (.CLK(clknet_4_3_0_wb_clk_i),
    .D(_0140_),
    .Q(\simon0.seq[19][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3358_ (.CLK(clknet_4_1_0_wb_clk_i),
    .D(_0141_),
    .Q(\simon0.seq[25][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3359_ (.CLK(clknet_4_1_0_wb_clk_i),
    .D(_0142_),
    .Q(\simon0.seq[25][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3360_ (.CLK(clknet_4_1_0_wb_clk_i),
    .D(_0143_),
    .Q(\simon0.seq[24][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3361_ (.CLK(clknet_4_1_0_wb_clk_i),
    .D(_0144_),
    .Q(\simon0.seq[24][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3362_ (.CLK(clknet_4_4_0_wb_clk_i),
    .D(_0145_),
    .Q(\simon0.seq[23][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3363_ (.CLK(clknet_4_4_0_wb_clk_i),
    .D(_0146_),
    .Q(\simon0.seq[23][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3364_ (.CLK(clknet_4_1_0_wb_clk_i),
    .D(_0147_),
    .Q(\simon0.seq[26][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3365_ (.CLK(clknet_4_1_0_wb_clk_i),
    .D(_0148_),
    .Q(\simon0.seq[26][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3366_ (.CLK(clknet_4_7_0_wb_clk_i),
    .D(_0149_),
    .Q(\simon0.seq[28][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3367_ (.CLK(clknet_4_7_0_wb_clk_i),
    .D(_0150_),
    .Q(\simon0.seq[28][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3368_ (.CLK(clknet_4_0_0_wb_clk_i),
    .D(_0151_),
    .Q(\simon0.seq[1][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3369_ (.CLK(clknet_4_0_0_wb_clk_i),
    .D(_0152_),
    .Q(\simon0.seq[1][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3370_ (.CLK(clknet_4_1_0_wb_clk_i),
    .D(_0153_),
    .Q(\simon0.seq[27][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3371_ (.CLK(clknet_4_1_0_wb_clk_i),
    .D(_0154_),
    .Q(\simon0.seq[27][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3372_ (.CLK(clknet_4_1_0_wb_clk_i),
    .D(_0155_),
    .Q(\simon0.seq[2][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3373_ (.CLK(clknet_4_1_0_wb_clk_i),
    .D(_0156_),
    .Q(\simon0.seq[2][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3374_ (.CLK(clknet_4_4_0_wb_clk_i),
    .D(_0157_),
    .Q(\simon0.seq[9][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3375_ (.CLK(clknet_4_4_0_wb_clk_i),
    .D(_0158_),
    .Q(\simon0.seq[9][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3376_ (.CLK(clknet_4_3_0_wb_clk_i),
    .D(_0159_),
    .Q(\simon0.seq[18][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3377_ (.CLK(clknet_4_3_0_wb_clk_i),
    .D(_0160_),
    .Q(\simon0.seq[18][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3378_ (.CLK(clknet_4_5_0_wb_clk_i),
    .D(_0161_),
    .Q(\simon0.seq[31][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3379_ (.CLK(clknet_4_5_0_wb_clk_i),
    .D(_0162_),
    .Q(\simon0.seq[31][1] ));
 sky130_fd_sc_hd__dfxtp_4 _3380_ (.CLK(clknet_4_6_0_wb_clk_i),
    .D(_0163_),
    .Q(_0000_));
 sky130_fd_sc_hd__dfxtp_2 _3381_ (.CLK(clknet_4_3_0_wb_clk_i),
    .D(_0164_),
    .Q(_0001_));
 sky130_fd_sc_hd__dfxtp_1 _3382_ (.CLK(clknet_4_6_0_wb_clk_i),
    .D(_0165_),
    .Q(_0002_));
 sky130_fd_sc_hd__dfxtp_1 _3383_ (.CLK(clknet_4_6_0_wb_clk_i),
    .D(_0166_),
    .Q(_0003_));
 sky130_fd_sc_hd__dfxtp_1 _3384_ (.CLK(clknet_4_2_0_wb_clk_i),
    .D(_0167_),
    .Q(_0004_));
 sky130_fd_sc_hd__dfxtp_1 _3385_ (.CLK(clknet_4_4_0_wb_clk_i),
    .D(_0168_),
    .Q(\simon0.seq[21][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3386_ (.CLK(clknet_4_4_0_wb_clk_i),
    .D(_0169_),
    .Q(\simon0.seq[21][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3387_ (.CLK(clknet_4_2_0_wb_clk_i),
    .D(_0170_),
    .Q(\simon0.seq[17][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3388_ (.CLK(clknet_4_2_0_wb_clk_i),
    .D(_0171_),
    .Q(\simon0.seq[17][1] ));
 sky130_fd_sc_hd__conb_1 _3493__25 (.LO(net25));
 sky130_fd_sc_hd__conb_1 _3494__26 (.LO(net26));
 sky130_fd_sc_hd__conb_1 _3495__27 (.LO(net27));
 sky130_fd_sc_hd__conb_1 _3496__28 (.LO(net28));
 sky130_fd_sc_hd__conb_1 _3497__29 (.LO(net29));
 sky130_fd_sc_hd__conb_1 _3498__30 (.LO(net30));
 sky130_fd_sc_hd__conb_1 _3499__31 (.LO(net31));
 sky130_fd_sc_hd__conb_1 _3500__32 (.LO(net32));
 sky130_fd_sc_hd__conb_1 _3501__33 (.LO(net33));
 sky130_fd_sc_hd__conb_1 _3502__34 (.LO(net34));
 sky130_fd_sc_hd__conb_1 _3503__35 (.LO(net35));
 sky130_fd_sc_hd__conb_1 _3504__36 (.LO(net36));
 sky130_fd_sc_hd__conb_1 _3505__37 (.LO(net37));
 sky130_fd_sc_hd__conb_1 _3506__38 (.LO(net38));
 sky130_fd_sc_hd__conb_1 _3507__39 (.LO(net39));
 sky130_fd_sc_hd__conb_1 _3508__40 (.LO(net40));
 sky130_fd_sc_hd__conb_1 _3509__41 (.LO(net41));
 sky130_fd_sc_hd__conb_1 _3510__42 (.LO(net42));
 sky130_fd_sc_hd__conb_1 _3511__43 (.LO(net43));
 sky130_fd_sc_hd__conb_1 _3512__44 (.LO(net44));
 sky130_fd_sc_hd__conb_1 _3513__45 (.LO(net45));
 sky130_fd_sc_hd__conb_1 _3514__46 (.LO(net46));
 sky130_fd_sc_hd__conb_1 _3515__47 (.LO(net47));
 sky130_fd_sc_hd__conb_1 _3516__48 (.LO(net48));
 sky130_fd_sc_hd__conb_1 _3517__49 (.LO(net49));
 sky130_fd_sc_hd__conb_1 _3518__50 (.LO(net50));
 sky130_fd_sc_hd__conb_1 _3519__51 (.LO(net51));
 sky130_fd_sc_hd__conb_1 _3520__52 (.LO(net52));
 sky130_fd_sc_hd__conb_1 _3521__53 (.LO(net53));
 sky130_fd_sc_hd__conb_1 _3522__54 (.LO(net54));
 sky130_fd_sc_hd__conb_1 _3523__55 (.LO(net55));
 sky130_fd_sc_hd__conb_1 _3524__56 (.LO(net56));
 sky130_fd_sc_hd__conb_1 _3525__57 (.LO(net57));
 sky130_fd_sc_hd__conb_1 _3526__58 (.LO(net58));
 sky130_fd_sc_hd__conb_1 _3527__59 (.LO(net59));
 sky130_fd_sc_hd__conb_1 _3528__60 (.LO(net60));
 sky130_fd_sc_hd__conb_1 _3529__61 (.LO(net61));
 sky130_fd_sc_hd__conb_1 _3530__62 (.LO(net62));
 sky130_fd_sc_hd__conb_1 _3531__63 (.LO(net63));
 sky130_fd_sc_hd__conb_1 _3532__64 (.LO(net64));
 sky130_fd_sc_hd__conb_1 _3533__65 (.LO(net65));
 sky130_fd_sc_hd__conb_1 _3534__66 (.LO(net66));
 sky130_fd_sc_hd__conb_1 _3535__67 (.LO(net67));
 sky130_fd_sc_hd__conb_1 _3541__68 (.LO(net68));
 sky130_fd_sc_hd__conb_1 _3542__69 (.LO(net69));
 sky130_fd_sc_hd__conb_1 _3543__70 (.LO(net70));
 sky130_fd_sc_hd__conb_1 _3544__71 (.LO(net71));
 sky130_fd_sc_hd__conb_1 _3545__72 (.LO(net72));
 sky130_fd_sc_hd__conb_1 _3546__73 (.LO(net73));
 sky130_fd_sc_hd__conb_1 _3547__74 (.LO(net74));
 sky130_fd_sc_hd__conb_1 _3548__75 (.LO(net75));
 sky130_fd_sc_hd__conb_1 _3549__76 (.LO(net76));
 sky130_fd_sc_hd__conb_1 _3550__77 (.LO(net77));
 sky130_fd_sc_hd__conb_1 _3551__78 (.LO(net78));
 sky130_fd_sc_hd__conb_1 _3552__79 (.LO(net79));
 sky130_fd_sc_hd__conb_1 _3553__80 (.LO(net80));
 sky130_fd_sc_hd__conb_1 _3554__81 (.LO(net81));
 sky130_fd_sc_hd__conb_1 _3555__82 (.LO(net82));
 sky130_fd_sc_hd__conb_1 _3556__83 (.LO(net83));
 sky130_fd_sc_hd__conb_1 _3557__84 (.LO(net84));
 sky130_fd_sc_hd__conb_1 _3558__85 (.LO(net85));
 sky130_fd_sc_hd__conb_1 _3559__86 (.LO(net86));
 sky130_fd_sc_hd__conb_1 _3560__87 (.LO(net87));
 sky130_fd_sc_hd__conb_1 _3561__88 (.LO(net88));
 sky130_fd_sc_hd__conb_1 _3562__89 (.LO(net89));
 sky130_fd_sc_hd__conb_1 _3563__90 (.LO(net90));
 sky130_fd_sc_hd__conb_1 _3564__91 (.LO(net91));
 sky130_fd_sc_hd__conb_1 _3565__92 (.LO(net92));
 sky130_fd_sc_hd__conb_1 _3566__93 (.LO(net93));
 sky130_fd_sc_hd__conb_1 _3567__94 (.LO(net94));
 sky130_fd_sc_hd__conb_1 _3568__95 (.LO(net95));
 sky130_fd_sc_hd__conb_1 _3569__96 (.LO(net96));
 sky130_fd_sc_hd__conb_1 _3570__97 (.LO(net97));
 sky130_fd_sc_hd__conb_1 _3571__98 (.LO(net98));
 sky130_fd_sc_hd__conb_1 _3572__99 (.LO(net99));
 sky130_fd_sc_hd__conb_1 _3573__100 (.LO(net100));
 sky130_fd_sc_hd__conb_1 _3574__101 (.LO(net101));
 sky130_fd_sc_hd__conb_1 _3575__102 (.LO(net102));
 sky130_fd_sc_hd__conb_1 _3576__103 (.LO(net103));
 sky130_fd_sc_hd__conb_1 _3577__104 (.LO(net104));
 sky130_fd_sc_hd__conb_1 _3578__105 (.LO(net105));
 sky130_fd_sc_hd__conb_1 _3579__106 (.LO(net106));
 sky130_fd_sc_hd__conb_1 _3580__107 (.LO(net107));
 sky130_fd_sc_hd__conb_1 _3581__108 (.LO(net108));
 sky130_fd_sc_hd__conb_1 _3582__109 (.LO(net109));
 sky130_fd_sc_hd__conb_1 _3583__110 (.LO(net110));
 sky130_fd_sc_hd__conb_1 _3584__111 (.LO(net111));
 sky130_fd_sc_hd__conb_1 _3585__112 (.LO(net112));
 sky130_fd_sc_hd__conb_1 _3586__113 (.LO(net113));
 sky130_fd_sc_hd__conb_1 _3587__114 (.LO(net114));
 sky130_fd_sc_hd__conb_1 _3588__115 (.LO(net115));
 sky130_fd_sc_hd__conb_1 _3589__116 (.LO(net116));
 sky130_fd_sc_hd__conb_1 _3590__117 (.LO(net117));
 sky130_fd_sc_hd__conb_1 _3591__118 (.LO(net118));
 sky130_fd_sc_hd__conb_1 _3592__119 (.LO(net119));
 sky130_fd_sc_hd__conb_1 _3593__120 (.LO(net120));
 sky130_fd_sc_hd__conb_1 _3594__121 (.LO(net121));
 sky130_fd_sc_hd__conb_1 _3595__122 (.LO(net122));
 sky130_fd_sc_hd__conb_1 _3596__123 (.LO(net123));
 sky130_fd_sc_hd__conb_1 _3597__124 (.LO(net124));
 sky130_fd_sc_hd__conb_1 _3598__125 (.LO(net125));
 sky130_fd_sc_hd__conb_1 _3599__126 (.LO(net126));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_wb_clk_i (.A(wb_clk_i),
    .X(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__ebufn_8 _3492_ (.A(net24),
    .TE_B(_1454_),
    .Z(la1_data_out[0]));
 sky130_fd_sc_hd__ebufn_8 _3493_ (.A(net25),
    .TE_B(_1455_),
    .Z(la1_data_out[1]));
 sky130_fd_sc_hd__ebufn_8 _3494_ (.A(net26),
    .TE_B(_1456_),
    .Z(la1_data_out[2]));
 sky130_fd_sc_hd__ebufn_8 _3495_ (.A(net27),
    .TE_B(_1457_),
    .Z(la1_data_out[3]));
 sky130_fd_sc_hd__ebufn_8 _3496_ (.A(net28),
    .TE_B(_1458_),
    .Z(la1_data_out[4]));
 sky130_fd_sc_hd__ebufn_8 _3497_ (.A(net29),
    .TE_B(_1459_),
    .Z(la1_data_out[5]));
 sky130_fd_sc_hd__ebufn_8 _3498_ (.A(net30),
    .TE_B(_1460_),
    .Z(la1_data_out[6]));
 sky130_fd_sc_hd__ebufn_8 _3499_ (.A(net31),
    .TE_B(_1461_),
    .Z(la1_data_out[7]));
 sky130_fd_sc_hd__ebufn_8 _3500_ (.A(net32),
    .TE_B(_1462_),
    .Z(la1_data_out[8]));
 sky130_fd_sc_hd__ebufn_8 _3501_ (.A(net33),
    .TE_B(_1463_),
    .Z(la1_data_out[9]));
 sky130_fd_sc_hd__ebufn_8 _3502_ (.A(net34),
    .TE_B(_1464_),
    .Z(la1_data_out[10]));
 sky130_fd_sc_hd__ebufn_8 _3503_ (.A(net35),
    .TE_B(_1465_),
    .Z(la1_data_out[11]));
 sky130_fd_sc_hd__ebufn_8 _3504_ (.A(net36),
    .TE_B(_1466_),
    .Z(la1_data_out[12]));
 sky130_fd_sc_hd__ebufn_8 _3505_ (.A(net37),
    .TE_B(_1467_),
    .Z(la1_data_out[13]));
 sky130_fd_sc_hd__ebufn_8 _3506_ (.A(net38),
    .TE_B(_1468_),
    .Z(la1_data_out[14]));
 sky130_fd_sc_hd__ebufn_8 _3507_ (.A(net39),
    .TE_B(_1469_),
    .Z(la1_data_out[15]));
 sky130_fd_sc_hd__ebufn_8 _3508_ (.A(net40),
    .TE_B(_1470_),
    .Z(la1_data_out[16]));
 sky130_fd_sc_hd__ebufn_8 _3509_ (.A(net41),
    .TE_B(_1471_),
    .Z(la1_data_out[17]));
 sky130_fd_sc_hd__ebufn_8 _3510_ (.A(net42),
    .TE_B(_1472_),
    .Z(la1_data_out[18]));
 sky130_fd_sc_hd__ebufn_8 _3511_ (.A(net43),
    .TE_B(_1473_),
    .Z(la1_data_out[19]));
 sky130_fd_sc_hd__ebufn_8 _3512_ (.A(net44),
    .TE_B(_1474_),
    .Z(la1_data_out[20]));
 sky130_fd_sc_hd__ebufn_8 _3513_ (.A(net45),
    .TE_B(_1475_),
    .Z(la1_data_out[21]));
 sky130_fd_sc_hd__ebufn_8 _3514_ (.A(net46),
    .TE_B(_1476_),
    .Z(la1_data_out[22]));
 sky130_fd_sc_hd__ebufn_8 _3515_ (.A(net47),
    .TE_B(_1477_),
    .Z(la1_data_out[23]));
 sky130_fd_sc_hd__ebufn_8 _3516_ (.A(net48),
    .TE_B(_1478_),
    .Z(la1_data_out[24]));
 sky130_fd_sc_hd__ebufn_8 _3517_ (.A(net49),
    .TE_B(_1479_),
    .Z(la1_data_out[25]));
 sky130_fd_sc_hd__ebufn_8 _3518_ (.A(net50),
    .TE_B(_1480_),
    .Z(la1_data_out[26]));
 sky130_fd_sc_hd__ebufn_8 _3519_ (.A(net51),
    .TE_B(_1481_),
    .Z(la1_data_out[27]));
 sky130_fd_sc_hd__ebufn_8 _3520_ (.A(net52),
    .TE_B(_1482_),
    .Z(la1_data_out[28]));
 sky130_fd_sc_hd__ebufn_8 _3521_ (.A(net53),
    .TE_B(_1483_),
    .Z(la1_data_out[29]));
 sky130_fd_sc_hd__ebufn_8 _3522_ (.A(net54),
    .TE_B(_1484_),
    .Z(la1_data_out[30]));
 sky130_fd_sc_hd__ebufn_8 _3523_ (.A(net55),
    .TE_B(_1485_),
    .Z(la1_data_out[31]));
 sky130_fd_sc_hd__ebufn_8 _3524_ (.A(net56),
    .TE_B(_1486_),
    .Z(io_out[0]));
 sky130_fd_sc_hd__ebufn_8 _3525_ (.A(net57),
    .TE_B(_1487_),
    .Z(io_out[1]));
 sky130_fd_sc_hd__ebufn_8 _3526_ (.A(net58),
    .TE_B(_1488_),
    .Z(io_out[2]));
 sky130_fd_sc_hd__ebufn_8 _3527_ (.A(net59),
    .TE_B(_1489_),
    .Z(io_out[3]));
 sky130_fd_sc_hd__ebufn_8 _3528_ (.A(net60),
    .TE_B(_1490_),
    .Z(io_out[4]));
 sky130_fd_sc_hd__ebufn_8 _3529_ (.A(net61),
    .TE_B(_1491_),
    .Z(io_out[5]));
 sky130_fd_sc_hd__ebufn_8 _3530_ (.A(net62),
    .TE_B(_1492_),
    .Z(io_out[6]));
 sky130_fd_sc_hd__ebufn_8 _3531_ (.A(net63),
    .TE_B(_1493_),
    .Z(io_out[7]));
 sky130_fd_sc_hd__ebufn_8 _3532_ (.A(net64),
    .TE_B(_1494_),
    .Z(io_out[8]));
 sky130_fd_sc_hd__ebufn_8 _3533_ (.A(net65),
    .TE_B(_1495_),
    .Z(io_out[9]));
 sky130_fd_sc_hd__ebufn_8 _3534_ (.A(net66),
    .TE_B(_1496_),
    .Z(io_out[10]));
 sky130_fd_sc_hd__ebufn_8 _3535_ (.A(net67),
    .TE_B(_1497_),
    .Z(io_out[11]));
 sky130_fd_sc_hd__ebufn_8 _3536_ (.A(\simon0.led[0] ),
    .TE_B(_1498_),
    .Z(io_out[12]));
 sky130_fd_sc_hd__ebufn_8 _3537_ (.A(\simon0.led[1] ),
    .TE_B(_1499_),
    .Z(io_out[13]));
 sky130_fd_sc_hd__ebufn_8 _3538_ (.A(\simon0.led[2] ),
    .TE_B(_1500_),
    .Z(io_out[14]));
 sky130_fd_sc_hd__ebufn_8 _3539_ (.A(\simon0.led[3] ),
    .TE_B(_1501_),
    .Z(io_out[15]));
 sky130_fd_sc_hd__ebufn_8 _3540_ (.A(\simon0.play1.sound ),
    .TE_B(_1502_),
    .Z(io_out[16]));
 sky130_fd_sc_hd__ebufn_8 _3541_ (.A(net68),
    .TE_B(_1503_),
    .Z(io_out[17]));
 sky130_fd_sc_hd__ebufn_8 _3542_ (.A(net69),
    .TE_B(_1504_),
    .Z(io_out[18]));
 sky130_fd_sc_hd__ebufn_8 _3543_ (.A(net70),
    .TE_B(_1505_),
    .Z(io_out[19]));
 sky130_fd_sc_hd__ebufn_8 _3544_ (.A(net71),
    .TE_B(_1506_),
    .Z(io_out[20]));
 sky130_fd_sc_hd__ebufn_8 _3545_ (.A(net72),
    .TE_B(_1507_),
    .Z(io_out[21]));
 sky130_fd_sc_hd__ebufn_8 _3546_ (.A(net73),
    .TE_B(_1508_),
    .Z(io_out[22]));
 sky130_fd_sc_hd__ebufn_8 _3547_ (.A(net74),
    .TE_B(_1509_),
    .Z(io_out[23]));
 sky130_fd_sc_hd__ebufn_8 _3548_ (.A(net75),
    .TE_B(_1510_),
    .Z(io_out[24]));
 sky130_fd_sc_hd__ebufn_8 _3549_ (.A(net76),
    .TE_B(_1511_),
    .Z(io_out[25]));
 sky130_fd_sc_hd__ebufn_8 _3550_ (.A(net77),
    .TE_B(_1512_),
    .Z(io_out[26]));
 sky130_fd_sc_hd__ebufn_8 _3551_ (.A(net78),
    .TE_B(_1513_),
    .Z(io_out[27]));
 sky130_fd_sc_hd__ebufn_8 _3552_ (.A(net79),
    .TE_B(_1514_),
    .Z(io_out[28]));
 sky130_fd_sc_hd__ebufn_8 _3553_ (.A(net80),
    .TE_B(_1515_),
    .Z(io_out[29]));
 sky130_fd_sc_hd__ebufn_8 _3554_ (.A(net81),
    .TE_B(_1516_),
    .Z(io_out[30]));
 sky130_fd_sc_hd__ebufn_8 _3555_ (.A(net82),
    .TE_B(_1517_),
    .Z(io_out[31]));
 sky130_fd_sc_hd__ebufn_8 _3556_ (.A(net83),
    .TE_B(_1518_),
    .Z(io_out[32]));
 sky130_fd_sc_hd__ebufn_8 _3557_ (.A(net84),
    .TE_B(_1519_),
    .Z(io_out[33]));
 sky130_fd_sc_hd__ebufn_8 _3558_ (.A(net85),
    .TE_B(_1520_),
    .Z(io_out[34]));
 sky130_fd_sc_hd__ebufn_8 _3559_ (.A(net86),
    .TE_B(_1521_),
    .Z(io_out[35]));
 sky130_fd_sc_hd__ebufn_8 _3560_ (.A(net87),
    .TE_B(_1522_),
    .Z(io_out[36]));
 sky130_fd_sc_hd__ebufn_8 _3561_ (.A(net88),
    .TE_B(_1523_),
    .Z(io_out[37]));
 sky130_fd_sc_hd__ebufn_8 _3562_ (.A(net89),
    .TE_B(_1524_),
    .Z(io_oeb[0]));
 sky130_fd_sc_hd__ebufn_8 _3563_ (.A(net90),
    .TE_B(_1525_),
    .Z(io_oeb[1]));
 sky130_fd_sc_hd__ebufn_8 _3564_ (.A(net91),
    .TE_B(_1526_),
    .Z(io_oeb[2]));
 sky130_fd_sc_hd__ebufn_8 _3565_ (.A(net92),
    .TE_B(_1527_),
    .Z(io_oeb[3]));
 sky130_fd_sc_hd__ebufn_8 _3566_ (.A(net93),
    .TE_B(_1528_),
    .Z(io_oeb[4]));
 sky130_fd_sc_hd__ebufn_8 _3567_ (.A(net94),
    .TE_B(_1529_),
    .Z(io_oeb[5]));
 sky130_fd_sc_hd__ebufn_8 _3568_ (.A(net95),
    .TE_B(_1530_),
    .Z(io_oeb[6]));
 sky130_fd_sc_hd__ebufn_8 _3569_ (.A(net96),
    .TE_B(_1531_),
    .Z(io_oeb[7]));
 sky130_fd_sc_hd__ebufn_8 _3570_ (.A(net97),
    .TE_B(_1532_),
    .Z(io_oeb[8]));
 sky130_fd_sc_hd__ebufn_8 _3571_ (.A(net98),
    .TE_B(_1533_),
    .Z(io_oeb[9]));
 sky130_fd_sc_hd__ebufn_8 _3572_ (.A(net99),
    .TE_B(_1534_),
    .Z(io_oeb[10]));
 sky130_fd_sc_hd__ebufn_8 _3573_ (.A(net100),
    .TE_B(_1535_),
    .Z(io_oeb[11]));
 sky130_fd_sc_hd__ebufn_8 _3574_ (.A(net101),
    .TE_B(_1536_),
    .Z(io_oeb[12]));
 sky130_fd_sc_hd__ebufn_8 _3575_ (.A(net102),
    .TE_B(_1537_),
    .Z(io_oeb[13]));
 sky130_fd_sc_hd__ebufn_8 _3576_ (.A(net103),
    .TE_B(_1538_),
    .Z(io_oeb[14]));
 sky130_fd_sc_hd__ebufn_8 _3577_ (.A(net104),
    .TE_B(_1539_),
    .Z(io_oeb[15]));
 sky130_fd_sc_hd__ebufn_8 _3578_ (.A(net105),
    .TE_B(_1540_),
    .Z(io_oeb[16]));
 sky130_fd_sc_hd__ebufn_8 _3579_ (.A(net106),
    .TE_B(_1541_),
    .Z(io_oeb[17]));
 sky130_fd_sc_hd__ebufn_8 _3580_ (.A(net107),
    .TE_B(_1542_),
    .Z(io_oeb[18]));
 sky130_fd_sc_hd__ebufn_8 _3581_ (.A(net108),
    .TE_B(_1543_),
    .Z(io_oeb[19]));
 sky130_fd_sc_hd__ebufn_8 _3582_ (.A(net109),
    .TE_B(_1544_),
    .Z(io_oeb[20]));
 sky130_fd_sc_hd__ebufn_8 _3583_ (.A(net110),
    .TE_B(_1545_),
    .Z(io_oeb[21]));
 sky130_fd_sc_hd__ebufn_8 _3584_ (.A(net111),
    .TE_B(_1546_),
    .Z(io_oeb[22]));
 sky130_fd_sc_hd__ebufn_8 _3585_ (.A(net112),
    .TE_B(_1547_),
    .Z(io_oeb[23]));
 sky130_fd_sc_hd__ebufn_8 _3586_ (.A(net113),
    .TE_B(_1548_),
    .Z(io_oeb[24]));
 sky130_fd_sc_hd__ebufn_8 _3587_ (.A(net114),
    .TE_B(_1549_),
    .Z(io_oeb[25]));
 sky130_fd_sc_hd__ebufn_8 _3588_ (.A(net115),
    .TE_B(_1550_),
    .Z(io_oeb[26]));
 sky130_fd_sc_hd__ebufn_8 _3589_ (.A(net116),
    .TE_B(_1551_),
    .Z(io_oeb[27]));
 sky130_fd_sc_hd__ebufn_8 _3590_ (.A(net117),
    .TE_B(_1552_),
    .Z(io_oeb[28]));
 sky130_fd_sc_hd__ebufn_8 _3591_ (.A(net118),
    .TE_B(_1553_),
    .Z(io_oeb[29]));
 sky130_fd_sc_hd__ebufn_8 _3592_ (.A(net119),
    .TE_B(_1554_),
    .Z(io_oeb[30]));
 sky130_fd_sc_hd__ebufn_8 _3593_ (.A(net120),
    .TE_B(_1555_),
    .Z(io_oeb[31]));
 sky130_fd_sc_hd__ebufn_8 _3594_ (.A(net121),
    .TE_B(_1556_),
    .Z(io_oeb[32]));
 sky130_fd_sc_hd__ebufn_8 _3595_ (.A(net122),
    .TE_B(_1557_),
    .Z(io_oeb[33]));
 sky130_fd_sc_hd__ebufn_8 _3596_ (.A(net123),
    .TE_B(_1558_),
    .Z(io_oeb[34]));
 sky130_fd_sc_hd__ebufn_8 _3597_ (.A(net124),
    .TE_B(_1559_),
    .Z(io_oeb[35]));
 sky130_fd_sc_hd__ebufn_8 _3598_ (.A(net125),
    .TE_B(_1560_),
    .Z(io_oeb[36]));
 sky130_fd_sc_hd__ebufn_8 _3599_ (.A(net126),
    .TE_B(_1561_),
    .Z(io_oeb[37]));
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__decap_3 PHY_92 ();
 sky130_fd_sc_hd__decap_3 PHY_93 ();
 sky130_fd_sc_hd__decap_3 PHY_94 ();
 sky130_fd_sc_hd__decap_3 PHY_95 ();
 sky130_fd_sc_hd__decap_3 PHY_96 ();
 sky130_fd_sc_hd__decap_3 PHY_97 ();
 sky130_fd_sc_hd__decap_3 PHY_98 ();
 sky130_fd_sc_hd__decap_3 PHY_99 ();
 sky130_fd_sc_hd__decap_3 PHY_100 ();
 sky130_fd_sc_hd__decap_3 PHY_101 ();
 sky130_fd_sc_hd__decap_3 PHY_102 ();
 sky130_fd_sc_hd__decap_3 PHY_103 ();
 sky130_fd_sc_hd__decap_3 PHY_104 ();
 sky130_fd_sc_hd__decap_3 PHY_105 ();
 sky130_fd_sc_hd__decap_3 PHY_106 ();
 sky130_fd_sc_hd__decap_3 PHY_107 ();
 sky130_fd_sc_hd__decap_3 PHY_108 ();
 sky130_fd_sc_hd__decap_3 PHY_109 ();
 sky130_fd_sc_hd__decap_3 PHY_110 ();
 sky130_fd_sc_hd__decap_3 PHY_111 ();
 sky130_fd_sc_hd__decap_3 PHY_112 ();
 sky130_fd_sc_hd__decap_3 PHY_113 ();
 sky130_fd_sc_hd__decap_3 PHY_114 ();
 sky130_fd_sc_hd__decap_3 PHY_115 ();
 sky130_fd_sc_hd__decap_3 PHY_116 ();
 sky130_fd_sc_hd__decap_3 PHY_117 ();
 sky130_fd_sc_hd__decap_3 PHY_118 ();
 sky130_fd_sc_hd__decap_3 PHY_119 ();
 sky130_fd_sc_hd__decap_3 PHY_120 ();
 sky130_fd_sc_hd__decap_3 PHY_121 ();
 sky130_fd_sc_hd__decap_3 PHY_122 ();
 sky130_fd_sc_hd__decap_3 PHY_123 ();
 sky130_fd_sc_hd__decap_3 PHY_124 ();
 sky130_fd_sc_hd__decap_3 PHY_125 ();
 sky130_fd_sc_hd__decap_3 PHY_126 ();
 sky130_fd_sc_hd__decap_3 PHY_127 ();
 sky130_fd_sc_hd__decap_3 PHY_128 ();
 sky130_fd_sc_hd__decap_3 PHY_129 ();
 sky130_fd_sc_hd__decap_3 PHY_130 ();
 sky130_fd_sc_hd__decap_3 PHY_131 ();
 sky130_fd_sc_hd__decap_3 PHY_132 ();
 sky130_fd_sc_hd__decap_3 PHY_133 ();
 sky130_fd_sc_hd__decap_3 PHY_134 ();
 sky130_fd_sc_hd__decap_3 PHY_135 ();
 sky130_fd_sc_hd__decap_3 PHY_136 ();
 sky130_fd_sc_hd__decap_3 PHY_137 ();
 sky130_fd_sc_hd__decap_3 PHY_138 ();
 sky130_fd_sc_hd__decap_3 PHY_139 ();
 sky130_fd_sc_hd__decap_3 PHY_140 ();
 sky130_fd_sc_hd__decap_3 PHY_141 ();
 sky130_fd_sc_hd__decap_3 PHY_142 ();
 sky130_fd_sc_hd__decap_3 PHY_143 ();
 sky130_fd_sc_hd__decap_3 PHY_144 ();
 sky130_fd_sc_hd__decap_3 PHY_145 ();
 sky130_fd_sc_hd__decap_3 PHY_146 ();
 sky130_fd_sc_hd__decap_3 PHY_147 ();
 sky130_fd_sc_hd__decap_3 PHY_148 ();
 sky130_fd_sc_hd__decap_3 PHY_149 ();
 sky130_fd_sc_hd__decap_3 PHY_150 ();
 sky130_fd_sc_hd__decap_3 PHY_151 ();
 sky130_fd_sc_hd__decap_3 PHY_152 ();
 sky130_fd_sc_hd__decap_3 PHY_153 ();
 sky130_fd_sc_hd__decap_3 PHY_154 ();
 sky130_fd_sc_hd__decap_3 PHY_155 ();
 sky130_fd_sc_hd__decap_3 PHY_156 ();
 sky130_fd_sc_hd__decap_3 PHY_157 ();
 sky130_fd_sc_hd__decap_3 PHY_158 ();
 sky130_fd_sc_hd__decap_3 PHY_159 ();
 sky130_fd_sc_hd__decap_3 PHY_160 ();
 sky130_fd_sc_hd__decap_3 PHY_161 ();
 sky130_fd_sc_hd__decap_3 PHY_162 ();
 sky130_fd_sc_hd__decap_3 PHY_163 ();
 sky130_fd_sc_hd__decap_3 PHY_164 ();
 sky130_fd_sc_hd__decap_3 PHY_165 ();
 sky130_fd_sc_hd__decap_3 PHY_166 ();
 sky130_fd_sc_hd__decap_3 PHY_167 ();
 sky130_fd_sc_hd__decap_3 PHY_168 ();
 sky130_fd_sc_hd__decap_3 PHY_169 ();
 sky130_fd_sc_hd__decap_3 PHY_170 ();
 sky130_fd_sc_hd__decap_3 PHY_171 ();
 sky130_fd_sc_hd__decap_3 PHY_172 ();
 sky130_fd_sc_hd__decap_3 PHY_173 ();
 sky130_fd_sc_hd__decap_3 PHY_174 ();
 sky130_fd_sc_hd__decap_3 PHY_175 ();
 sky130_fd_sc_hd__decap_3 PHY_176 ();
 sky130_fd_sc_hd__decap_3 PHY_177 ();
 sky130_fd_sc_hd__decap_3 PHY_178 ();
 sky130_fd_sc_hd__decap_3 PHY_179 ();
 sky130_fd_sc_hd__decap_3 PHY_180 ();
 sky130_fd_sc_hd__decap_3 PHY_181 ();
 sky130_fd_sc_hd__decap_3 PHY_182 ();
 sky130_fd_sc_hd__decap_3 PHY_183 ();
 sky130_fd_sc_hd__decap_3 PHY_184 ();
 sky130_fd_sc_hd__decap_3 PHY_185 ();
 sky130_fd_sc_hd__decap_3 PHY_186 ();
 sky130_fd_sc_hd__decap_3 PHY_187 ();
 sky130_fd_sc_hd__decap_3 PHY_188 ();
 sky130_fd_sc_hd__decap_3 PHY_189 ();
 sky130_fd_sc_hd__decap_3 PHY_190 ();
 sky130_fd_sc_hd__decap_3 PHY_191 ();
 sky130_fd_sc_hd__decap_3 PHY_192 ();
 sky130_fd_sc_hd__decap_3 PHY_193 ();
 sky130_fd_sc_hd__decap_3 PHY_194 ();
 sky130_fd_sc_hd__decap_3 PHY_195 ();
 sky130_fd_sc_hd__decap_3 PHY_196 ();
 sky130_fd_sc_hd__decap_3 PHY_197 ();
 sky130_fd_sc_hd__decap_3 PHY_198 ();
 sky130_fd_sc_hd__decap_3 PHY_199 ();
 sky130_fd_sc_hd__decap_3 PHY_200 ();
 sky130_fd_sc_hd__decap_3 PHY_201 ();
 sky130_fd_sc_hd__decap_3 PHY_202 ();
 sky130_fd_sc_hd__decap_3 PHY_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1347 ();
 sky130_fd_sc_hd__clkbuf_1 input1 (.A(active),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_1 input2 (.A(io_in[10]),
    .X(net2));
 sky130_fd_sc_hd__buf_2 input3 (.A(io_in[11]),
    .X(net3));
 sky130_fd_sc_hd__buf_6 input4 (.A(io_in[17]),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_4 input5 (.A(io_in[18]),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_2 input6 (.A(io_in[8]),
    .X(net6));
 sky130_fd_sc_hd__buf_2 input7 (.A(io_in[9]),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_4 input8 (.A(la1_data_in[0]),
    .X(net8));
 sky130_fd_sc_hd__dlymetal6s2s_1 input9 (.A(la1_data_in[10]),
    .X(net9));
 sky130_fd_sc_hd__clkbuf_2 input10 (.A(la1_data_in[11]),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_4 input11 (.A(la1_data_in[12]),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_1 input12 (.A(la1_data_in[13]),
    .X(net12));
 sky130_fd_sc_hd__dlymetal6s2s_1 input13 (.A(la1_data_in[14]),
    .X(net13));
 sky130_fd_sc_hd__clkbuf_4 input14 (.A(la1_data_in[15]),
    .X(net14));
 sky130_fd_sc_hd__clkbuf_4 input15 (.A(la1_data_in[1]),
    .X(net15));
 sky130_fd_sc_hd__clkbuf_4 input16 (.A(la1_data_in[2]),
    .X(net16));
 sky130_fd_sc_hd__buf_2 input17 (.A(la1_data_in[3]),
    .X(net17));
 sky130_fd_sc_hd__buf_4 input18 (.A(la1_data_in[4]),
    .X(net18));
 sky130_fd_sc_hd__clkbuf_4 input19 (.A(la1_data_in[5]),
    .X(net19));
 sky130_fd_sc_hd__clkbuf_4 input20 (.A(la1_data_in[6]),
    .X(net20));
 sky130_fd_sc_hd__buf_2 input21 (.A(la1_data_in[7]),
    .X(net21));
 sky130_fd_sc_hd__clkbuf_4 input22 (.A(la1_data_in[8]),
    .X(net22));
 sky130_fd_sc_hd__buf_2 input23 (.A(la1_data_in[9]),
    .X(net23));
 sky130_fd_sc_hd__conb_1 _3492__24 (.LO(net24));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_0_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_4_0_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_1_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_4_1_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_2_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_4_2_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_3_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_4_3_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_4_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_4_4_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_5_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_4_5_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_6_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_4_6_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_7_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_4_7_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_8_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_4_8_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_9_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_4_9_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_10_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_4_10_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_11_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_4_11_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_12_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_4_12_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_13_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_4_13_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_14_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_4_14_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_15_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_4_15_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(\simon0.led[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2 (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA_3 (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA_4 (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA_5 (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA_6 (.DIODE(net11));
 sky130_fd_sc_hd__fill_2 FILLER_0_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_622 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_25 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_94 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_298 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_310 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_384 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_424 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_501 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_532 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_604 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_50 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_102 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_136 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_158 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_192 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_272 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_346 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_407 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_556 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_612 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_619 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_88 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_146 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_324 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_328 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_343 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_355 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_473 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_535 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_542 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_554 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_581 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_588 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_592 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_622 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_26 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_623 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_34 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_42 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_236 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_622 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_16 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_623 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_34 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_585 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_606 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_622 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_16 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_245 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_263 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_208 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_227 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_623 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_34 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_240 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_252 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_319 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_346 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_473 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_16 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_267 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_351 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_235 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_255 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_355 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_267 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_336 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_340 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_242 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_263 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_294 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_186 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_198 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_257 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_294 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_332 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_16 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_192 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_224 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_267 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_318 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_34 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_16 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_190 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_226 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_430 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_623 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_182 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_245 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_272 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_364 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_431 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_460 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_467 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_597 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_25 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_224 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_236 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_358 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_379 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_403 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_439 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_178 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_254 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_266 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_375 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_466 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_597 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_622 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_203 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_211 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_228 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_240 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_282 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_340 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_387 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_443 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_612 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_619 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_272 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_410 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_219 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_286 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_315 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_392 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_404 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_451 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_623 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_243 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_411 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_423 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_431 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_460 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_478 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_612 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_12 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_175 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_232 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_336 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_403 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_484 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_508 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_623 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_34 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_186 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_198 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_204 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_230 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_242 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_254 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_311 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_344 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_367 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_442 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_458 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_16 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_211 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_296 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_326 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_336 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_348 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_370 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_395 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_434 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_452 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_458 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_484 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_491 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_187 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_212 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_239 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_247 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_290 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_378 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_413 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_420 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_436 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_459 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_470 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_476 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_483 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_322 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_450 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_465 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_504 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_623 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_34 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_176 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_185 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_203 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_256 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_328 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_359 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_364 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_402 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_422 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_442 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_605 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_327 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_414 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_431 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_438 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_450 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_486 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_623 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_180 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_196 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_308 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_347 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_406 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_422 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_432 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_442 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_455 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_473 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_16 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_328 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_394 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_402 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_434 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_493 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_198 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_317 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_357 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_425 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_442 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_466 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_478 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_511 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_535 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_168 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_239 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_506 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_199 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_218 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_236 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_254 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_411 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_612 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_183 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_336 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_400 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_428 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_455 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_520 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_623 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_34 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_267 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_311 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_467 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_516 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_16 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_219 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_261 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_318 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_374 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_400 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_623 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_187 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_198 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_304 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_347 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_429 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_585 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_596 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_602 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_606 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_16 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_210 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_316 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_336 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_426 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_438 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_450 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_618 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_201 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_308 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_332 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_480 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_516 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_540 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_597 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_176 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_184 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_212 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_327 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_338 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_465 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_493 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_504 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_512 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_34 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_149 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_180 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_255 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_263 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_297 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_364 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_376 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_413 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_478 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_488 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_522 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_220 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_240 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_273 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_283 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_291 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_338 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_410 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_474 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_495 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_504 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_14 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_186 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_411 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_423 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_476 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_480 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_502 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_16 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_219 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_396 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_441 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_452 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_460 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_490 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_502 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_510 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_623 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_128 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_189 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_198 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_355 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_378 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_384 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_473 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_152 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_284 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_439 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_443 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_131 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_241 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_267 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_296 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_355 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_366 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_467 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_612 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_136 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_164 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_450 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_463 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_470 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_143 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_164 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_256 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_300 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_320 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_358 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_366 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_426 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_460 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_540 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_126 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_171 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_219 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_270 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_282 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_294 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_374 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_394 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_432 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_120 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_127 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_190 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_348 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_360 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_368 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_612 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_266 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_282 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_318 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_325 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_414 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_431 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_463 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_123 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_174 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_186 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_198 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_206 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_268 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_303 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_318 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_375 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_398 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_585 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_606 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_622 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_156 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_227 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_239 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_271 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_290 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_316 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_395 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_430 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_130 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_147 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_239 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_310 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_355 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_367 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_400 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_415 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_444 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_455 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_119 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_168 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_216 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_226 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_318 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_338 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_350 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_380 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_232 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_459 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_471 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_215 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_352 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_379 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_439 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_316 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_605 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_610 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_115 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_123 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_159 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_271 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_283 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_439 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_482 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_494 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_506 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_623 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_34 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_119 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_142 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_152 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_230 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_328 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_102 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_172 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_314 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_326 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_338 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_448 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_486 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_87 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_180 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_214 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_242 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_299 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_310 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_319 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_424 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_470 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_482 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_107 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_159 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_274 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_336 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_392 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_450 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_123 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_154 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_174 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_299 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_355 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_367 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_398 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_416 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_424 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_457 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_114 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_168 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_387 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_396 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_460 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_499 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_243 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_255 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_303 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_346 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_460 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_470 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_511 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_535 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_612 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_96 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_152 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_180 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_383 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_395 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_442 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_450 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_458 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_106 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_201 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_236 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_252 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_314 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_428 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_456 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_116 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_236 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_336 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_340 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_387 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_395 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_403 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_451 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_459 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_470 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_493 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_500 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_512 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_94 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_106 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_143 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_186 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_312 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_324 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_359 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_370 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_426 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_478 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_502 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_511 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_536 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_597 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_182 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_282 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_342 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_432 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_450 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_454 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_493 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_551 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_563 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_609 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_144 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_201 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_357 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_487 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_498 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_513 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_612 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_171 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_178 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_331 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_343 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_428 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_435 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_482 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_499 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_511 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_540 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_549 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_305 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_422 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_471 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_494 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_524 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_536 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_622 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_224 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_372 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_451 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_493 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_531 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_542 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_551 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_563 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_176 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_188 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_200 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_243 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_270 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_286 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_298 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_346 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_368 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_380 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_432 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_455 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_471 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_478 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_534 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_605 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_610 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_122 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_132 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_180 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_407 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_444 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_543 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_550 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_562 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_623 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_34 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_142 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_154 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_187 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_254 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_305 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_459 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_466 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_525 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_543 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_612 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_14 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_107 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_132 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_163 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_218 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_276 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_288 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_296 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_398 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_428 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_457 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_484 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_498 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_510 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_518 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_549 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_566 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_609 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_120 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_144 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_186 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_190 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_328 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_386 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_482 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_525 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_229 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_320 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_370 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_410 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_431 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_443 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_492 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_510 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_518 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_551 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_563 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_22 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_124 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_207 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_243 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_255 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_313 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_367 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_413 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_432 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_501 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_511 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_622 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_159 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_314 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_326 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_338 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_394 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_414 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_432 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_472 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_490 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_34 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_148 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_236 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_438 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_491 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_612 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_12 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_276 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_320 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_403 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_442 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_484 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_23 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_75 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_187 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_322 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_342 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_376 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_413 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_437 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_462 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_217 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_296 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_322 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_188 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_260 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_473 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_494 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_622 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_11 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_43 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_190 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_206 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_226 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_273 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_398 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_12 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_34 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_211 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_368 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_622 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_16 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_34 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_42 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_64 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_129 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_202 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_214 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_226 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_263 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_283 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_344 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_379 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_426 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_438 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_450 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_568 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_586 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_92 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_151 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_398 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_478 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_536 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_622 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_66 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_129 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_202 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_214 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_226 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_322 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_378 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_426 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_438 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_450 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_466 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_36 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_42 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_586 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_622 ();
endmodule

